-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : whiterabbit_gtpe2_channel_wrapper.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module whiterabbit_gtpe2_channel_wrapper (a GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

use work.wr_gtp_phy_pkg.all;

--***************************** Entity Declaration ****************************

entity whiterabbit_gtpe2_channel_wrapper is
generic
(
    -- Simulation attributes
    PLL0_FBDIV                     : integer := 4;
    PLL0_FBDIV_45                  : integer := 5;
    PLL0_REFCLK_DIV                : integer := 1;
    PLL1_FBDIV                     : integer := 4;
    PLL1_FBDIV_45                  : integer := 5;
    PLL1_REFCLK_DIV                : integer := 1;
    g_num_phys                     : integer := 1;
    EXAMPLE_SIMULATION             : integer  := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "true" to speed up sim reset
);
port
(
    GT_CHANNEL_SIG_i               : in   t_gtpe2_channel_in_array(g_num_phys-1 downto 0);
    GT_CHANNEL_SIG_o               : out  t_gtpe2_channel_out_array(g_num_phys-1 downto 0);
    -----------------------------COMMON PORTS-----------------------------------
    ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
    GTREFCLK0                      : in   std_logic;
    GTREFCLK1                      : in   std_logic;
    ----------------- Select the input reference clock to the CPLL -------------
    PLL0REFCLKSEL                  : in   std_logic_vector:="001";
    PLL1REFCLKSEL                  : in   std_logic_vector:="001";
    -------------------------- Common Block - PLL Ports ------------------------
    PLL0PD                         : in   std_logic:='0';
    PLL1PD                         : in   std_logic:='0';
    PLL0RESET                      : in   std_logic:='0';
    PLL1RESET                      : in   std_logic:='0';
    PLL0LOCK                       : out  std_logic;
    PLL1LOCK                       : out  std_logic;
    PLL0REFCLKLOST                 : out  std_logic;
    PLL1REFCLKLOST                 : out  std_logic;

    PLL0OUTCLK_OUT                 : out  std_logic;
    PLL0OUTREFCLK_OUT              : out  std_logic;
    PLL0LOCK_OUT                   : out  std_logic;
    PLL0LOCKDETCLK_IN              : in   std_logic;
    PLL0REFCLKLOST_OUT             : out  std_logic;
    PLL0RESET_IN                   : in   std_logic
);


end whiterabbit_gtpe2_channel_wrapper;
    
architecture RTL of whiterabbit_gtpe2_channel_wrapper is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "whiterabbit_gtpe2_channel_wrapper,gtwizard_v3_6_1,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i        :   std_logic;
    signal  tied_to_ground_vec_i    :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i           :   std_logic;

    signal  PLL0OUTCLK              :   std_logic;
    signal  PLL1OUTCLK              :   std_logic;
    signal  PLL0OUTREFCLK           :   std_logic;
    signal  PLL1OUTREFCLK           :   std_logic;
 
--*************************** Component Declarations **************************
component whiterabbit_gtpe2_channel_wrapper_gt
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "false";
    EXAMPLE_SIMULATION        : integer:= 0;  
    TXSYNC_OVRD_IN            : bit    := '0';
    TXSYNC_MULTILANE_IN       : bit    := '0'
);
port 
(
    ---------------------------- Channel - Reset   -----------------------------   
    RST_IN                                  : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    DRPADDR_IN                              : in   std_logic_vector(8 downto 0);
    DRPCLK_IN                               : in   std_logic;
    DRPDI_IN                                : in   std_logic_vector(15 downto 0);
    DRPDO_OUT                               : out  std_logic_vector(15 downto 0);
    DRPEN_IN                                : in   std_logic;
    DRPRDY_OUT                              : out  std_logic;
    DRPWE_IN                                : in   std_logic;
    DRP_BUSY_OUT                            : out  std_logic;
    ------------------------ GTPE2_CHANNEL Clocking Ports ----------------------
    RXSYSCLKSEL_IN                          : in   std_logic_vector(1 downto 0);
    TXSYSCLKSEL_IN                          : in   std_logic_vector(1 downto 0);
    PLL0CLK_IN                              : in   std_logic;
    PLL0REFCLK_IN                           : in   std_logic;
    PLL1CLK_IN                              : in   std_logic;
    PLL1REFCLK_IN                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    LOOPBACK_IN                             : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    RXUSERRDY_IN                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    EYESCANDATAERROR_OUT                    : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    RXDATA_OUT                              : out  std_logic_vector(31 downto 0);
    RXUSRCLK_IN                             : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    RXCHARISCOMMA_OUT                       : out  std_logic_vector(3 downto 0);
    RXCHARISK_OUT                           : out  std_logic_vector(3 downto 0);
    RXDISPERR_OUT                           : out  std_logic_vector(3 downto 0);
    RXNOTINTABLE_OUT                        : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GTPRXN_IN                               : in   std_logic;
    GTPRXP_IN                               : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    RXBYTEISALIGNED_OUT                     : out  std_logic;
    RXCOMMADET_OUT                          : out  std_logic;
    RXSLIDE_IN                              : in   std_logic;
    --------------------- Receive Ports - RX Equilizer Ports -------------------
    RXLPMHFHOLD_IN                          : in   std_logic;
    RXLPMLFHOLD_IN                          : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    RXOUTCLK_OUT                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GTRXRESET_IN                            : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    RXRESETDONE_OUT                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GTTXRESET_IN                            : in   std_logic;
    TXUSERRDY_IN                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    TXDATA_IN                               : in   std_logic_vector(31 downto 0);
    TXUSRCLK_IN                             : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    TXCHARISK_IN                            : in   std_logic_vector(3 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    GTPTXN_OUT                              : out  std_logic;
    GTPTXP_OUT                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    TXOUTCLK_OUT                            : out  std_logic;
    TXOUTCLKFABRIC_OUT                      : out  std_logic;
    TXOUTCLKPCS_OUT                         : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    TXRESETDONE_OUT                         : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    TXPRBSSEL_IN                            : in   std_logic_vector(2 downto 0)
);
end component;

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';

    --------------------------- GTPE2_COMMON -------------------------------
    gtpe2_common_0_i : GTPE2_COMMON
    generic map
    (
        -- Simulation attributes
        SIM_RESET_SPEEDUP               => WRAPPER_SIM_GTRESET_SPEEDUP,
        SIM_PLL0REFCLK_SEL              => ("001"),
        SIM_PLL1REFCLK_SEL              => ("001"),
        SIM_VERSION                     => ("1.0"),

        PLL0_FBDIV                      => PLL0_FBDIV,
        PLL0_FBDIV_45                   => PLL0_FBDIV_45,
        PLL0_REFCLK_DIV                 => PLL0_REFCLK_DIV,
        PLL1_FBDIV                      => PLL1_FBDIV,
        PLL1_FBDIV_45                   => PLL1_FBDIV_45,
        PLL1_REFCLK_DIV                 => PLL1_REFCLK_DIV,

       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                        =>     (x"0000000000050001"),
        COMMON_CFG                      =>     (x"00000000"),

       ----------------------------PLL Attributes----------------------------
        PLL0_CFG                        =>     (x"01F03DC"),
        PLL0_DMON_CFG                   =>     ('0'),
        PLL0_INIT_CFG                   =>     (x"00001E"),
        PLL0_LOCK_CFG                   =>     (x"1E8"),
        PLL1_CFG                        =>     (x"01F03DC"),
        PLL1_DMON_CFG                   =>     ('0'),
        PLL1_INIT_CFG                   =>     (x"00001E"),
        PLL1_LOCK_CFG                   =>     (x"1E8"),
        PLL_CLKOUT_CFG                  =>     (x"00"),

       ----------------------------Reserved Attributes----------------------------
        RSVD_ATTR0                      =>     (x"0000"),
        RSVD_ATTR1                      =>     (x"0000")
    )
    port map
    (
        DMONITOROUT                     =>      open,
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
        GTGREFCLK0                      =>      tied_to_ground_i,
        GTGREFCLK1                      =>      tied_to_ground_i,
        GTREFCLK0                       =>      GTREFCLK0,
        GTREFCLK1                       =>      GTREFCLK1,
        GTWESTREFCLK0                   =>      tied_to_ground_i,
        GTWESTREFCLK1                   =>      tied_to_ground_i,
        GTEASTREFCLK0                   =>      tied_to_ground_i,
        GTEASTREFCLK1                   =>      tied_to_ground_i,
        PLL0OUTCLK                      =>      PLL0OUTCLK_OUT,
        PLL1OUTCLK                      =>      PLL1OUTCLK,
        PLL0OUTREFCLK                   =>      PLL0OUTREFCLK_OUT,
        PLL1OUTREFCLK                   =>      PLL1OUTREFCLK,
        PLL0REFCLKSEL                   =>      PLL0REFCLKSEL,
        PLL1REFCLKSEL                   =>      PLL1REFCLKSEL,
        -------------------------- Common Block - PLL Ports ------------------------
        PLL0LOCKDETCLK                  =>      PLL0LOCKDETCLK_IN,
        PLL1LOCKDETCLK                  =>      tied_to_ground_i,
        PLL0LOCKEN                      =>      tied_to_vcc_i,
        PLL1LOCKEN                      =>      tied_to_vcc_i,
        PLL0PD                          =>      PLL0PD,
        PLL1PD                          =>      PLL1PD,
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "11111",
        RCALENB                         =>      tied_to_vcc_i,
        PLL0RESET                       =>      PLL0RESET_IN,
        PLL1RESET                       =>      PLL1RESET,
        PLL0FBCLKLOST                   =>      open,
        PLL1FBCLKLOST                   =>      open,
        PLL0LOCK                        =>      PLL0LOCK_OUT,
        PLL1LOCK                        =>      PLL1LOCK,
        PLL0REFCLKLOST                  =>      PLL0REFCLKLOST_OUT,
        PLL1REFCLKLOST                  =>      PLL1REFCLKLOST,
        ---------------------------- Common Block - Ports --------------------------
        BGRCALOVRDENB                   =>      tied_to_vcc_i,
        PLLRSVD1                        =>      "0000000000000000",
        PLLRSVD2                        =>      "00000",
        REFCLKOUTMONITOR0               =>      open,
        REFCLKOUTMONITOR1               =>      open,
        ------------------------ Common Block - RX AFE Ports -----------------------
        PMARSVDOUT                      =>      open,
        --------------------------------- QPLL Ports -------------------------------
        PMARSVD                         =>      "00000000"
    );

gen_GT_INTS: for i in 0 to g_num_phys-1 generate

    GT_INST : whiterabbit_gtpe2_channel_wrapper_gt
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        PLL0CLK_IN                      =>      PLL0OUTCLK,
        PLL0REFCLK_IN                   =>      PLL0OUTREFCLK,
        PLL1CLK_IN                      =>      PLL1OUTCLK,
        PLL1REFCLK_IN                   =>      PLL1OUTREFCLK,
        RST_IN                          =>      GT_CHANNEL_SIG_i(i).RST_IN,
        DRP_BUSY_OUT                    =>      GT_CHANNEL_SIG_o(i).DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT_CHANNEL_SIG_i(i).DRPADDR_IN,
        DRPCLK_IN                       =>      GT_CHANNEL_SIG_i(i).DRPCLK_IN,
        DRPDI_IN                        =>      GT_CHANNEL_SIG_i(i).DRPDI_IN,
        DRPDO_OUT                       =>      GT_CHANNEL_SIG_o(i).DRPDO_OUT,
        DRPEN_IN                        =>      GT_CHANNEL_SIG_i(i).DRPEN_IN,
        DRPRDY_OUT                      =>      GT_CHANNEL_SIG_o(i).DRPRDY_OUT,
        DRPWE_IN                        =>      GT_CHANNEL_SIG_i(i).DRPWE_IN,
        ------------------------ GTPE2_CHANNEL Clocking Ports ----------------------
        RXSYSCLKSEL_IN                  =>      GT_CHANNEL_SIG_i(i).RXSYSCLKSEL,
        TXSYSCLKSEL_IN                  =>      GT_CHANNEL_SIG_i(i).TXSYSCLKSEL,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT_CHANNEL_SIG_i(i).LOOPBACK,
        --------------------- RX Initialization and Reset Ports -------------------
        RXUSERRDY_IN                    =>      GT_CHANNEL_SIG_i(i).RXUSERRDY,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT_CHANNEL_SIG_o(i).EYESCANDATAERROR,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXDATA_OUT                      =>      GT_CHANNEL_SIG_o(i).RXDATA,
        RXUSRCLK_IN                     =>      GT_CHANNEL_SIG_i(i).RXUSRCLK,
        RXUSRCLK2_IN                    =>      GT_CHANNEL_SIG_i(i).RXUSRCLK2,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT_CHANNEL_SIG_o(i).RXCHARISCOMMA,
        RXCHARISK_OUT                   =>      GT_CHANNEL_SIG_o(i).RXCHARISK,
        RXDISPERR_OUT                   =>      GT_CHANNEL_SIG_o(i).RXDISPERR,
        RXNOTINTABLE_OUT                =>      GT_CHANNEL_SIG_o(i).RXNOTINTABLE,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTPRXN_IN                       =>      GT_CHANNEL_SIG_i(i).GTPRXN,
        GTPRXP_IN                       =>      GT_CHANNEL_SIG_i(i).GTPRXP,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT_CHANNEL_SIG_o(i).RXBYTEISALIGNED,
        RXCOMMADET_OUT                  =>      GT_CHANNEL_SIG_o(i).RXCOMMADET,
        RXSLIDE_IN                      =>      GT_CHANNEL_SIG_i(i).RXSLIDE,
        --------------------- Receive Ports - RX Equilizer Ports -------------------
        RXLPMHFHOLD_IN                  =>      GT_CHANNEL_SIG_i(i).RXLPMHFHOLD,
        RXLPMLFHOLD_IN                  =>      GT_CHANNEL_SIG_i(i).RXLPMLFHOLD,
        --------------- Receive Ports - RX Fabric Output Control Pors -------------
        RXOUTCLK_OUT                    =>      GT_CHANNEL_SIG_o(i).RXOUTCLK,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT_CHANNEL_SIG_i(i).GTRXRESET,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT_CHANNEL_SIG_o(i).RXRESETDONE,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT_CHANNEL_SIG_i(i).GTTXRESET,
        TXUSERRDY_IN                    =>      GT_CHANNEL_SIG_i(i).TXUSERRDY,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXDATA_IN                       =>      GT_CHANNEL_SIG_i(i).TXDATA,
        TXUSRCLK_IN                     =>      GT_CHANNEL_SIG_i(i).TXUSRCLK,
        TXUSRCLK2_IN                    =>      GT_CHANNEL_SIG_i(i).TXUSRCLK2,
        ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        TXCHARISK_IN                    =>      GT_CHANNEL_SIG_i(i).TXCHARISK,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        GTPTXN_OUT                      =>      GT_CHANNEL_SIG_o(i).GTPTXN,
        GTPTXP_OUT                      =>      GT_CHANNEL_SIG_o(i).GTPTXP,
        ----------- Transmit Ports - TX Fabric Clock Output Control ports ----------
        TXOUTCLK_OUT                    =>      GT_CHANNEL_SIG_o(i).TXOUTCLK,
        TXOUTCLKFABRIC_OUT              =>      GT_CHANNEL_SIG_o(i).TXOUTCLKFABRIC,
        TXOUTCLKPCS_OUT                 =>      GT_CHANNEL_SIG_o(i).TXOUTCLKPCS,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT_CHANNEL_SIG_o(i).TXRESETDONE,
        ------------------ Transmit Ports - pattern Generator Ports ---------------
        TXPRBSSEL_IN                    =>      GT_CHANNEL_SIG_i(i).TXPRBSSEL
    );
end generate gen_GT_INTS;

end RTL;
