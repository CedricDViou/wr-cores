// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "06/19/2019 10:23:20"

// 
// Device: Altera 10AX115S2F45I1SG Package FBGA1932
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module wr_arria10_e3p1_det_phy (
	reconfig_write,
	reconfig_read,
	reconfig_address,
	reconfig_writedata,
	reconfig_readdata,
	reconfig_waitrequest,
	reconfig_clk,
	reconfig_reset,
	rx_analogreset,
	rx_cal_busy,
	rx_cdr_refclk0,
	rx_clkout,
	rx_coreclkin,
	rx_datak,
	rx_digitalreset,
	rx_disperr,
	rx_errdetect,
	rx_is_lockedtodata,
	rx_is_lockedtoref,
	rx_parallel_data,
	rx_patterndetect,
	rx_runningdisp,
	rx_serial_data,
	rx_seriallpbken,
	rx_std_bitslipboundarysel,
	rx_std_wa_patternalign,
	rx_syncstatus,
	tx_analogreset,
	tx_cal_busy,
	tx_clkout,
	tx_coreclkin,
	tx_datak,
	tx_digitalreset,
	tx_parallel_data,
	tx_serial_clk0,
	tx_serial_data,
	unused_rx_parallel_data,
	unused_tx_parallel_data)/* synthesis synthesis_greybox=1 */;
input 	[0:0] reconfig_write;
input 	[0:0] reconfig_read;
input 	[9:0] reconfig_address;
input 	[31:0] reconfig_writedata;
output 	[31:0] reconfig_readdata;
output 	[0:0] reconfig_waitrequest;
input 	[0:0] reconfig_clk;
input 	[0:0] reconfig_reset;
input 	[0:0] rx_analogreset;
output 	[0:0] rx_cal_busy;
input 	rx_cdr_refclk0;
output 	[0:0] rx_clkout;
input 	[0:0] rx_coreclkin;
output 	rx_datak;
input 	[0:0] rx_digitalreset;
output 	rx_disperr;
output 	rx_errdetect;
output 	[0:0] rx_is_lockedtodata;
output 	[0:0] rx_is_lockedtoref;
output 	[7:0] rx_parallel_data;
output 	rx_patterndetect;
output 	rx_runningdisp;
input 	[0:0] rx_serial_data;
input 	[0:0] rx_seriallpbken;
output 	[4:0] rx_std_bitslipboundarysel;
input 	[0:0] rx_std_wa_patternalign;
output 	rx_syncstatus;
input 	[0:0] tx_analogreset;
output 	[0:0] tx_cal_busy;
output 	[0:0] tx_clkout;
input 	[0:0] tx_coreclkin;
input 	tx_datak;
input 	[0:0] tx_digitalreset;
input 	[7:0] tx_parallel_data;
input 	[0:0] tx_serial_clk0;
output 	[0:0] tx_serial_data;
output 	[113:0] unused_rx_parallel_data;
input 	[118:0] unused_tx_parallel_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[0] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[1] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[2] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[3] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[4] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[5] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[6] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[7] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[8] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[9] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[10] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[11] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[12] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[13] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[14] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[15] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[16] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[17] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[18] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[19] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[20] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[21] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[22] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[23] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[24] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[25] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[26] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[27] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[28] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[29] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[30] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[31] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[32] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[33] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[34] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[35] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[36] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[37] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[38] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[39] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[40] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[41] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[42] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[43] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[44] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[45] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[46] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[47] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[48] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[49] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[50] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[51] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[52] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[53] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[54] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[55] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[56] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[57] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[58] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[59] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[60] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[61] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[62] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[63] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[64] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[65] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[66] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[67] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[68] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[69] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[70] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[71] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[72] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[73] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[74] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[75] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[76] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[77] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[78] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[79] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[80] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[81] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[82] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[83] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[84] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[85] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[86] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[87] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[88] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[89] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[90] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[91] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[92] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[93] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[94] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[95] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[96] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[97] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[98] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[99] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[100] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[101] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[102] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[103] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[104] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[105] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[106] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[107] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[108] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[109] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[110] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[111] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[112] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[113] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[114] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[115] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[116] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[117] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[118] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[119] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[120] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[121] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[122] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[123] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[124] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[125] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[126] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[127] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|pld_cal_done[0] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[0] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[1] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[2] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[3] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[4] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[5] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[6] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[7] ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pma|w_pma_tx_buf_vop ;
wire \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_waitrequest[0]~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \reconfig_address[9]~input_o ;
wire \reconfig_writedata[8]~input_o ;
wire \reconfig_writedata[9]~input_o ;
wire \reconfig_writedata[10]~input_o ;
wire \reconfig_writedata[11]~input_o ;
wire \reconfig_writedata[12]~input_o ;
wire \reconfig_writedata[13]~input_o ;
wire \reconfig_writedata[14]~input_o ;
wire \reconfig_writedata[15]~input_o ;
wire \reconfig_writedata[16]~input_o ;
wire \reconfig_writedata[17]~input_o ;
wire \reconfig_writedata[18]~input_o ;
wire \reconfig_writedata[19]~input_o ;
wire \reconfig_writedata[20]~input_o ;
wire \reconfig_writedata[21]~input_o ;
wire \reconfig_writedata[22]~input_o ;
wire \reconfig_writedata[23]~input_o ;
wire \reconfig_writedata[24]~input_o ;
wire \reconfig_writedata[25]~input_o ;
wire \reconfig_writedata[26]~input_o ;
wire \reconfig_writedata[27]~input_o ;
wire \reconfig_writedata[28]~input_o ;
wire \reconfig_writedata[29]~input_o ;
wire \reconfig_writedata[30]~input_o ;
wire \reconfig_writedata[31]~input_o ;
wire \reconfig_read[0]~input_o ;
wire \tx_analogreset[0]~input_o ;
wire \rx_analogreset[0]~input_o ;
wire \rx_digitalreset[0]~input_o ;
wire \rx_std_wa_patternalign[0]~input_o ;
wire \rx_coreclkin[0]~input_o ;
wire \reconfig_clk[0]~input_o ;
wire \reconfig_write[0]~input_o ;
wire \reconfig_address[0]~input_o ;
wire \reconfig_address[1]~input_o ;
wire \reconfig_address[2]~input_o ;
wire \reconfig_address[3]~input_o ;
wire \reconfig_address[4]~input_o ;
wire \reconfig_address[5]~input_o ;
wire \reconfig_address[6]~input_o ;
wire \reconfig_address[7]~input_o ;
wire \reconfig_address[8]~input_o ;
wire \reconfig_writedata[0]~input_o ;
wire \reconfig_writedata[1]~input_o ;
wire \reconfig_writedata[2]~input_o ;
wire \reconfig_writedata[3]~input_o ;
wire \reconfig_writedata[4]~input_o ;
wire \reconfig_writedata[5]~input_o ;
wire \reconfig_writedata[6]~input_o ;
wire \reconfig_writedata[7]~input_o ;
wire \rx_seriallpbken[0]~input_o ;
wire \tx_digitalreset[0]~input_o ;
wire \tx_coreclkin[0]~input_o ;
wire \tx_parallel_data[0]~input_o ;
wire \tx_parallel_data[1]~input_o ;
wire \tx_parallel_data[2]~input_o ;
wire \tx_parallel_data[3]~input_o ;
wire \tx_parallel_data[4]~input_o ;
wire \tx_parallel_data[5]~input_o ;
wire \tx_parallel_data[6]~input_o ;
wire \tx_parallel_data[7]~input_o ;
wire \tx_datak~input_o ;
wire \unused_tx_parallel_data[0]~input_o ;
wire \unused_tx_parallel_data[1]~input_o ;
wire \unused_tx_parallel_data[2]~input_o ;
wire \unused_tx_parallel_data[3]~input_o ;
wire \unused_tx_parallel_data[4]~input_o ;
wire \unused_tx_parallel_data[5]~input_o ;
wire \unused_tx_parallel_data[6]~input_o ;
wire \unused_tx_parallel_data[7]~input_o ;
wire \unused_tx_parallel_data[8]~input_o ;
wire \unused_tx_parallel_data[9]~input_o ;
wire \unused_tx_parallel_data[10]~input_o ;
wire \unused_tx_parallel_data[11]~input_o ;
wire \unused_tx_parallel_data[12]~input_o ;
wire \unused_tx_parallel_data[13]~input_o ;
wire \unused_tx_parallel_data[14]~input_o ;
wire \unused_tx_parallel_data[15]~input_o ;
wire \unused_tx_parallel_data[16]~input_o ;
wire \unused_tx_parallel_data[17]~input_o ;
wire \unused_tx_parallel_data[18]~input_o ;
wire \unused_tx_parallel_data[19]~input_o ;
wire \unused_tx_parallel_data[20]~input_o ;
wire \unused_tx_parallel_data[21]~input_o ;
wire \unused_tx_parallel_data[22]~input_o ;
wire \unused_tx_parallel_data[23]~input_o ;
wire \unused_tx_parallel_data[24]~input_o ;
wire \unused_tx_parallel_data[25]~input_o ;
wire \unused_tx_parallel_data[26]~input_o ;
wire \unused_tx_parallel_data[27]~input_o ;
wire \unused_tx_parallel_data[28]~input_o ;
wire \unused_tx_parallel_data[29]~input_o ;
wire \unused_tx_parallel_data[30]~input_o ;
wire \unused_tx_parallel_data[31]~input_o ;
wire \unused_tx_parallel_data[32]~input_o ;
wire \unused_tx_parallel_data[33]~input_o ;
wire \unused_tx_parallel_data[34]~input_o ;
wire \unused_tx_parallel_data[35]~input_o ;
wire \unused_tx_parallel_data[36]~input_o ;
wire \unused_tx_parallel_data[37]~input_o ;
wire \unused_tx_parallel_data[38]~input_o ;
wire \unused_tx_parallel_data[39]~input_o ;
wire \unused_tx_parallel_data[40]~input_o ;
wire \unused_tx_parallel_data[41]~input_o ;
wire \unused_tx_parallel_data[42]~input_o ;
wire \unused_tx_parallel_data[43]~input_o ;
wire \unused_tx_parallel_data[44]~input_o ;
wire \unused_tx_parallel_data[45]~input_o ;
wire \unused_tx_parallel_data[46]~input_o ;
wire \unused_tx_parallel_data[47]~input_o ;
wire \unused_tx_parallel_data[48]~input_o ;
wire \unused_tx_parallel_data[49]~input_o ;
wire \unused_tx_parallel_data[50]~input_o ;
wire \unused_tx_parallel_data[51]~input_o ;
wire \unused_tx_parallel_data[52]~input_o ;
wire \unused_tx_parallel_data[53]~input_o ;
wire \unused_tx_parallel_data[54]~input_o ;
wire \unused_tx_parallel_data[55]~input_o ;
wire \unused_tx_parallel_data[56]~input_o ;
wire \unused_tx_parallel_data[57]~input_o ;
wire \unused_tx_parallel_data[58]~input_o ;
wire \unused_tx_parallel_data[59]~input_o ;
wire \unused_tx_parallel_data[60]~input_o ;
wire \unused_tx_parallel_data[61]~input_o ;
wire \unused_tx_parallel_data[62]~input_o ;
wire \unused_tx_parallel_data[63]~input_o ;
wire \unused_tx_parallel_data[64]~input_o ;
wire \unused_tx_parallel_data[65]~input_o ;
wire \unused_tx_parallel_data[66]~input_o ;
wire \unused_tx_parallel_data[67]~input_o ;
wire \unused_tx_parallel_data[68]~input_o ;
wire \unused_tx_parallel_data[69]~input_o ;
wire \unused_tx_parallel_data[70]~input_o ;
wire \unused_tx_parallel_data[71]~input_o ;
wire \unused_tx_parallel_data[72]~input_o ;
wire \unused_tx_parallel_data[73]~input_o ;
wire \unused_tx_parallel_data[74]~input_o ;
wire \unused_tx_parallel_data[75]~input_o ;
wire \unused_tx_parallel_data[76]~input_o ;
wire \unused_tx_parallel_data[77]~input_o ;
wire \unused_tx_parallel_data[78]~input_o ;
wire \unused_tx_parallel_data[79]~input_o ;
wire \unused_tx_parallel_data[80]~input_o ;
wire \unused_tx_parallel_data[81]~input_o ;
wire \unused_tx_parallel_data[82]~input_o ;
wire \unused_tx_parallel_data[83]~input_o ;
wire \unused_tx_parallel_data[84]~input_o ;
wire \unused_tx_parallel_data[85]~input_o ;
wire \unused_tx_parallel_data[86]~input_o ;
wire \unused_tx_parallel_data[87]~input_o ;
wire \unused_tx_parallel_data[88]~input_o ;
wire \unused_tx_parallel_data[89]~input_o ;
wire \unused_tx_parallel_data[90]~input_o ;
wire \unused_tx_parallel_data[91]~input_o ;
wire \unused_tx_parallel_data[92]~input_o ;
wire \unused_tx_parallel_data[93]~input_o ;
wire \unused_tx_parallel_data[94]~input_o ;
wire \unused_tx_parallel_data[95]~input_o ;
wire \unused_tx_parallel_data[96]~input_o ;
wire \unused_tx_parallel_data[97]~input_o ;
wire \unused_tx_parallel_data[98]~input_o ;
wire \unused_tx_parallel_data[99]~input_o ;
wire \unused_tx_parallel_data[100]~input_o ;
wire \unused_tx_parallel_data[101]~input_o ;
wire \unused_tx_parallel_data[102]~input_o ;
wire \unused_tx_parallel_data[103]~input_o ;
wire \unused_tx_parallel_data[104]~input_o ;
wire \unused_tx_parallel_data[105]~input_o ;
wire \unused_tx_parallel_data[106]~input_o ;
wire \unused_tx_parallel_data[107]~input_o ;
wire \unused_tx_parallel_data[108]~input_o ;
wire \unused_tx_parallel_data[109]~input_o ;
wire \unused_tx_parallel_data[110]~input_o ;
wire \unused_tx_parallel_data[111]~input_o ;
wire \unused_tx_parallel_data[112]~input_o ;
wire \unused_tx_parallel_data[113]~input_o ;
wire \unused_tx_parallel_data[114]~input_o ;
wire \unused_tx_parallel_data[115]~input_o ;
wire \unused_tx_parallel_data[116]~input_o ;
wire \unused_tx_parallel_data[117]~input_o ;
wire \unused_tx_parallel_data[118]~input_o ;
wire \rx_serial_data[0]~input_o ;
wire \tx_serial_clk0[0]~input_o ;
wire \rx_cdr_refclk0~input_o ;
wire \reconfig_reset[0]~input_o ;


wr_arria10_e3p1_det_phy_wr_arria10_e3p1_det_phy_altera_xcvr_native_a10_181_iwfuxyq xcvr_native_a10_0(
	.w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out ),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0] ),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1] ),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2] ),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3] ),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_0(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[0] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_1(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[1] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_2(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[2] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_3(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[3] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_4(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[4] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_5(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[5] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_6(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[6] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_7(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[7] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_8(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[8] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_9(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[9] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_10(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[10] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_11(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[11] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_12(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[12] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_13(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[13] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_14(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[14] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_15(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[15] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_16(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[16] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_17(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[17] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_18(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[18] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_19(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[19] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_20(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[20] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_21(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[21] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_22(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[22] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_23(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[23] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_24(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[24] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_25(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[25] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_26(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[26] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_27(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[27] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_28(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[28] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_29(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[29] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_30(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[30] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_31(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[31] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_32(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[32] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_33(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[33] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_34(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[34] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_35(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[35] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_36(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[36] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_37(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[37] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_38(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[38] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_39(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[39] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_40(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[40] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_41(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[41] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_42(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[42] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_43(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[43] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_44(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[44] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_45(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[45] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_46(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[46] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_47(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[47] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_48(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[48] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_49(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[49] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_50(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[50] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_51(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[51] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_52(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[52] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_53(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[53] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_54(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[54] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_55(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[55] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_56(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[56] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_57(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[57] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_58(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[58] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_59(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[59] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_60(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[60] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_61(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[61] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_62(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[62] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_63(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[63] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_64(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[64] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_65(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[65] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_66(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[66] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_67(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[67] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_68(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[68] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_69(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[69] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_70(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[70] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_71(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[71] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_72(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[72] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_73(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[73] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_74(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[74] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_75(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[75] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_76(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[76] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_77(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[77] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_78(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[78] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_79(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[79] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_80(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[80] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_81(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[81] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_82(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[82] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_83(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[83] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_84(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[84] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_85(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[85] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_86(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[86] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_87(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[87] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_88(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[88] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_89(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[89] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_90(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[90] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_91(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[91] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_92(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[92] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_93(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[93] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_94(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[94] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_95(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[95] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_96(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[96] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_97(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[97] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_98(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[98] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_99(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[99] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_100(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[100] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_101(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[101] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_102(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[102] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_103(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[103] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_104(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[104] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_105(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[105] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_106(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[106] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_107(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[107] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_108(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[108] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_109(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[109] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_110(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[110] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_111(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[111] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_112(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[112] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_113(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[113] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_114(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[114] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_115(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[115] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_116(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[116] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_117(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[117] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_118(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[118] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_119(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[119] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_120(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[120] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_121(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[121] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_122(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[122] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_123(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[123] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_124(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[124] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_125(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[125] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_126(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[126] ),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_127(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[127] ),
	.pld_cal_done_0(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|pld_cal_done[0] ),
	.avmm_readdata_0(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[0] ),
	.avmm_readdata_1(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[1] ),
	.avmm_readdata_2(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[2] ),
	.avmm_readdata_3(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[3] ),
	.avmm_readdata_4(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[4] ),
	.avmm_readdata_5(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[5] ),
	.avmm_readdata_6(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[6] ),
	.avmm_readdata_7(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[7] ),
	.w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock ),
	.w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock ),
	.tx_clkout({\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out }),
	.tx_serial_data({\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pma|w_pma_tx_buf_vop }),
	.avmm_waitrequest_0(\xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_waitrequest[0]~0_combout ),
	.reset_out_stage_0(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0]~q ),
	.reset_out_stage_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1]~q ),
	.reconfig_read_0(\reconfig_read[0]~input_o ),
	.rx_digitalreset_0(\rx_digitalreset[0]~input_o ),
	.rx_std_wa_patternalign_0(\rx_std_wa_patternalign[0]~input_o ),
	.rx_coreclkin_0(\rx_coreclkin[0]~input_o ),
	.reconfig_clk_0(\reconfig_clk[0]~input_o ),
	.reconfig_write_0(\reconfig_write[0]~input_o ),
	.reconfig_address_0(\reconfig_address[0]~input_o ),
	.reconfig_address_1(\reconfig_address[1]~input_o ),
	.reconfig_address_2(\reconfig_address[2]~input_o ),
	.reconfig_address_3(\reconfig_address[3]~input_o ),
	.reconfig_address_4(\reconfig_address[4]~input_o ),
	.reconfig_address_5(\reconfig_address[5]~input_o ),
	.reconfig_address_6(\reconfig_address[6]~input_o ),
	.reconfig_address_7(\reconfig_address[7]~input_o ),
	.reconfig_address_8(\reconfig_address[8]~input_o ),
	.reconfig_writedata_0(\reconfig_writedata[0]~input_o ),
	.reconfig_writedata_1(\reconfig_writedata[1]~input_o ),
	.reconfig_writedata_2(\reconfig_writedata[2]~input_o ),
	.reconfig_writedata_3(\reconfig_writedata[3]~input_o ),
	.reconfig_writedata_4(\reconfig_writedata[4]~input_o ),
	.reconfig_writedata_5(\reconfig_writedata[5]~input_o ),
	.reconfig_writedata_6(\reconfig_writedata[6]~input_o ),
	.reconfig_writedata_7(\reconfig_writedata[7]~input_o ),
	.rx_seriallpbken_0(\rx_seriallpbken[0]~input_o ),
	.tx_digitalreset_0(\tx_digitalreset[0]~input_o ),
	.tx_coreclkin_0(\tx_coreclkin[0]~input_o ),
	.tx_parallel_data_0(\tx_parallel_data[0]~input_o ),
	.tx_parallel_data_1(\tx_parallel_data[1]~input_o ),
	.tx_parallel_data_2(\tx_parallel_data[2]~input_o ),
	.tx_parallel_data_3(\tx_parallel_data[3]~input_o ),
	.tx_parallel_data_4(\tx_parallel_data[4]~input_o ),
	.tx_parallel_data_5(\tx_parallel_data[5]~input_o ),
	.tx_parallel_data_6(\tx_parallel_data[6]~input_o ),
	.tx_parallel_data_7(\tx_parallel_data[7]~input_o ),
	.tx_datak(\tx_datak~input_o ),
	.unused_tx_parallel_data_0(\unused_tx_parallel_data[0]~input_o ),
	.unused_tx_parallel_data_1(\unused_tx_parallel_data[1]~input_o ),
	.unused_tx_parallel_data_2(\unused_tx_parallel_data[2]~input_o ),
	.unused_tx_parallel_data_3(\unused_tx_parallel_data[3]~input_o ),
	.unused_tx_parallel_data_4(\unused_tx_parallel_data[4]~input_o ),
	.unused_tx_parallel_data_5(\unused_tx_parallel_data[5]~input_o ),
	.unused_tx_parallel_data_6(\unused_tx_parallel_data[6]~input_o ),
	.unused_tx_parallel_data_7(\unused_tx_parallel_data[7]~input_o ),
	.unused_tx_parallel_data_8(\unused_tx_parallel_data[8]~input_o ),
	.unused_tx_parallel_data_9(\unused_tx_parallel_data[9]~input_o ),
	.unused_tx_parallel_data_10(\unused_tx_parallel_data[10]~input_o ),
	.unused_tx_parallel_data_11(\unused_tx_parallel_data[11]~input_o ),
	.unused_tx_parallel_data_12(\unused_tx_parallel_data[12]~input_o ),
	.unused_tx_parallel_data_13(\unused_tx_parallel_data[13]~input_o ),
	.unused_tx_parallel_data_14(\unused_tx_parallel_data[14]~input_o ),
	.unused_tx_parallel_data_15(\unused_tx_parallel_data[15]~input_o ),
	.unused_tx_parallel_data_16(\unused_tx_parallel_data[16]~input_o ),
	.unused_tx_parallel_data_17(\unused_tx_parallel_data[17]~input_o ),
	.unused_tx_parallel_data_18(\unused_tx_parallel_data[18]~input_o ),
	.unused_tx_parallel_data_19(\unused_tx_parallel_data[19]~input_o ),
	.unused_tx_parallel_data_20(\unused_tx_parallel_data[20]~input_o ),
	.unused_tx_parallel_data_21(\unused_tx_parallel_data[21]~input_o ),
	.unused_tx_parallel_data_22(\unused_tx_parallel_data[22]~input_o ),
	.unused_tx_parallel_data_23(\unused_tx_parallel_data[23]~input_o ),
	.unused_tx_parallel_data_24(\unused_tx_parallel_data[24]~input_o ),
	.unused_tx_parallel_data_25(\unused_tx_parallel_data[25]~input_o ),
	.unused_tx_parallel_data_26(\unused_tx_parallel_data[26]~input_o ),
	.unused_tx_parallel_data_27(\unused_tx_parallel_data[27]~input_o ),
	.unused_tx_parallel_data_28(\unused_tx_parallel_data[28]~input_o ),
	.unused_tx_parallel_data_29(\unused_tx_parallel_data[29]~input_o ),
	.unused_tx_parallel_data_30(\unused_tx_parallel_data[30]~input_o ),
	.unused_tx_parallel_data_31(\unused_tx_parallel_data[31]~input_o ),
	.unused_tx_parallel_data_32(\unused_tx_parallel_data[32]~input_o ),
	.unused_tx_parallel_data_33(\unused_tx_parallel_data[33]~input_o ),
	.unused_tx_parallel_data_34(\unused_tx_parallel_data[34]~input_o ),
	.unused_tx_parallel_data_35(\unused_tx_parallel_data[35]~input_o ),
	.unused_tx_parallel_data_36(\unused_tx_parallel_data[36]~input_o ),
	.unused_tx_parallel_data_37(\unused_tx_parallel_data[37]~input_o ),
	.unused_tx_parallel_data_38(\unused_tx_parallel_data[38]~input_o ),
	.unused_tx_parallel_data_39(\unused_tx_parallel_data[39]~input_o ),
	.unused_tx_parallel_data_40(\unused_tx_parallel_data[40]~input_o ),
	.unused_tx_parallel_data_41(\unused_tx_parallel_data[41]~input_o ),
	.unused_tx_parallel_data_42(\unused_tx_parallel_data[42]~input_o ),
	.unused_tx_parallel_data_43(\unused_tx_parallel_data[43]~input_o ),
	.unused_tx_parallel_data_44(\unused_tx_parallel_data[44]~input_o ),
	.unused_tx_parallel_data_45(\unused_tx_parallel_data[45]~input_o ),
	.unused_tx_parallel_data_46(\unused_tx_parallel_data[46]~input_o ),
	.unused_tx_parallel_data_47(\unused_tx_parallel_data[47]~input_o ),
	.unused_tx_parallel_data_48(\unused_tx_parallel_data[48]~input_o ),
	.unused_tx_parallel_data_49(\unused_tx_parallel_data[49]~input_o ),
	.unused_tx_parallel_data_50(\unused_tx_parallel_data[50]~input_o ),
	.unused_tx_parallel_data_51(\unused_tx_parallel_data[51]~input_o ),
	.unused_tx_parallel_data_52(\unused_tx_parallel_data[52]~input_o ),
	.unused_tx_parallel_data_53(\unused_tx_parallel_data[53]~input_o ),
	.unused_tx_parallel_data_54(\unused_tx_parallel_data[54]~input_o ),
	.unused_tx_parallel_data_55(\unused_tx_parallel_data[55]~input_o ),
	.unused_tx_parallel_data_56(\unused_tx_parallel_data[56]~input_o ),
	.unused_tx_parallel_data_57(\unused_tx_parallel_data[57]~input_o ),
	.unused_tx_parallel_data_58(\unused_tx_parallel_data[58]~input_o ),
	.unused_tx_parallel_data_59(\unused_tx_parallel_data[59]~input_o ),
	.unused_tx_parallel_data_60(\unused_tx_parallel_data[60]~input_o ),
	.unused_tx_parallel_data_61(\unused_tx_parallel_data[61]~input_o ),
	.unused_tx_parallel_data_62(\unused_tx_parallel_data[62]~input_o ),
	.unused_tx_parallel_data_63(\unused_tx_parallel_data[63]~input_o ),
	.unused_tx_parallel_data_64(\unused_tx_parallel_data[64]~input_o ),
	.unused_tx_parallel_data_65(\unused_tx_parallel_data[65]~input_o ),
	.unused_tx_parallel_data_66(\unused_tx_parallel_data[66]~input_o ),
	.unused_tx_parallel_data_67(\unused_tx_parallel_data[67]~input_o ),
	.unused_tx_parallel_data_68(\unused_tx_parallel_data[68]~input_o ),
	.unused_tx_parallel_data_69(\unused_tx_parallel_data[69]~input_o ),
	.unused_tx_parallel_data_70(\unused_tx_parallel_data[70]~input_o ),
	.unused_tx_parallel_data_71(\unused_tx_parallel_data[71]~input_o ),
	.unused_tx_parallel_data_72(\unused_tx_parallel_data[72]~input_o ),
	.unused_tx_parallel_data_73(\unused_tx_parallel_data[73]~input_o ),
	.unused_tx_parallel_data_74(\unused_tx_parallel_data[74]~input_o ),
	.unused_tx_parallel_data_75(\unused_tx_parallel_data[75]~input_o ),
	.unused_tx_parallel_data_76(\unused_tx_parallel_data[76]~input_o ),
	.unused_tx_parallel_data_77(\unused_tx_parallel_data[77]~input_o ),
	.unused_tx_parallel_data_78(\unused_tx_parallel_data[78]~input_o ),
	.unused_tx_parallel_data_79(\unused_tx_parallel_data[79]~input_o ),
	.unused_tx_parallel_data_80(\unused_tx_parallel_data[80]~input_o ),
	.unused_tx_parallel_data_81(\unused_tx_parallel_data[81]~input_o ),
	.unused_tx_parallel_data_82(\unused_tx_parallel_data[82]~input_o ),
	.unused_tx_parallel_data_83(\unused_tx_parallel_data[83]~input_o ),
	.unused_tx_parallel_data_84(\unused_tx_parallel_data[84]~input_o ),
	.unused_tx_parallel_data_85(\unused_tx_parallel_data[85]~input_o ),
	.unused_tx_parallel_data_86(\unused_tx_parallel_data[86]~input_o ),
	.unused_tx_parallel_data_87(\unused_tx_parallel_data[87]~input_o ),
	.unused_tx_parallel_data_88(\unused_tx_parallel_data[88]~input_o ),
	.unused_tx_parallel_data_89(\unused_tx_parallel_data[89]~input_o ),
	.unused_tx_parallel_data_90(\unused_tx_parallel_data[90]~input_o ),
	.unused_tx_parallel_data_91(\unused_tx_parallel_data[91]~input_o ),
	.unused_tx_parallel_data_92(\unused_tx_parallel_data[92]~input_o ),
	.unused_tx_parallel_data_93(\unused_tx_parallel_data[93]~input_o ),
	.unused_tx_parallel_data_94(\unused_tx_parallel_data[94]~input_o ),
	.unused_tx_parallel_data_95(\unused_tx_parallel_data[95]~input_o ),
	.unused_tx_parallel_data_96(\unused_tx_parallel_data[96]~input_o ),
	.unused_tx_parallel_data_97(\unused_tx_parallel_data[97]~input_o ),
	.unused_tx_parallel_data_98(\unused_tx_parallel_data[98]~input_o ),
	.unused_tx_parallel_data_99(\unused_tx_parallel_data[99]~input_o ),
	.unused_tx_parallel_data_100(\unused_tx_parallel_data[100]~input_o ),
	.unused_tx_parallel_data_101(\unused_tx_parallel_data[101]~input_o ),
	.unused_tx_parallel_data_102(\unused_tx_parallel_data[102]~input_o ),
	.unused_tx_parallel_data_103(\unused_tx_parallel_data[103]~input_o ),
	.unused_tx_parallel_data_104(\unused_tx_parallel_data[104]~input_o ),
	.unused_tx_parallel_data_105(\unused_tx_parallel_data[105]~input_o ),
	.unused_tx_parallel_data_106(\unused_tx_parallel_data[106]~input_o ),
	.unused_tx_parallel_data_107(\unused_tx_parallel_data[107]~input_o ),
	.unused_tx_parallel_data_108(\unused_tx_parallel_data[108]~input_o ),
	.unused_tx_parallel_data_109(\unused_tx_parallel_data[109]~input_o ),
	.unused_tx_parallel_data_110(\unused_tx_parallel_data[110]~input_o ),
	.unused_tx_parallel_data_111(\unused_tx_parallel_data[111]~input_o ),
	.unused_tx_parallel_data_112(\unused_tx_parallel_data[112]~input_o ),
	.unused_tx_parallel_data_113(\unused_tx_parallel_data[113]~input_o ),
	.unused_tx_parallel_data_114(\unused_tx_parallel_data[114]~input_o ),
	.unused_tx_parallel_data_115(\unused_tx_parallel_data[115]~input_o ),
	.unused_tx_parallel_data_116(\unused_tx_parallel_data[116]~input_o ),
	.unused_tx_parallel_data_117(\unused_tx_parallel_data[117]~input_o ),
	.unused_tx_parallel_data_118(\unused_tx_parallel_data[118]~input_o ),
	.rx_serial_data_0(\rx_serial_data[0]~input_o ),
	.tx_serial_clk0_0(\tx_serial_clk0[0]~input_o ),
	.rx_cdr_refclk0(\rx_cdr_refclk0~input_o ),
	.reconfig_reset_0(\reconfig_reset[0]~input_o ));

twentynm_oscillator \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS (
	.oscena(!\auto_hub|~GND~combout ),
	.clkout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.clkout1());

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_stage[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0] .power_up = "low";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0 .lut_mask = 64'h5FFF5FFFF5FFF5FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2] .power_up = "low";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[1] .power_up = "low";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~0 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1 .lut_mask = 64'hDFFDFDDFFDDFDFFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~1 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2 .lut_mask = 64'hFF7DFF7DFF7DFF7D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~2 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\tx_analogreset[0]~input_o ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[0].sync_r[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(\rx_analogreset[0]~input_o ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[2]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0] (
	.clk(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|ALTERA_INSERTED_INTOSC_FOR_TRS~clkout ),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_n_generator|resync_chains[0].sync_r[0] .power_up = "low";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_match~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_counter~4 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|Equal0~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_req_synchronizers|resync_chains[1].sync_r[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|sched_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:without_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|a10xcvrfabric|altera_reset_sequencer|reset_out_reg[1]~1 .shared_arith = "off";

twentynm_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

assign \reconfig_read[0]~input_o  = reconfig_read[0];

assign \tx_analogreset[0]~input_o  = tx_analogreset[0];

assign \rx_analogreset[0]~input_o  = rx_analogreset[0];

assign \rx_digitalreset[0]~input_o  = rx_digitalreset[0];

assign \rx_std_wa_patternalign[0]~input_o  = rx_std_wa_patternalign[0];

assign \rx_coreclkin[0]~input_o  = rx_coreclkin[0];

assign \reconfig_clk[0]~input_o  = reconfig_clk[0];

assign \reconfig_write[0]~input_o  = reconfig_write[0];

assign \reconfig_address[0]~input_o  = reconfig_address[0];

assign \reconfig_address[1]~input_o  = reconfig_address[1];

assign \reconfig_address[2]~input_o  = reconfig_address[2];

assign \reconfig_address[3]~input_o  = reconfig_address[3];

assign \reconfig_address[4]~input_o  = reconfig_address[4];

assign \reconfig_address[5]~input_o  = reconfig_address[5];

assign \reconfig_address[6]~input_o  = reconfig_address[6];

assign \reconfig_address[7]~input_o  = reconfig_address[7];

assign \reconfig_address[8]~input_o  = reconfig_address[8];

assign \reconfig_writedata[0]~input_o  = reconfig_writedata[0];

assign \reconfig_writedata[1]~input_o  = reconfig_writedata[1];

assign \reconfig_writedata[2]~input_o  = reconfig_writedata[2];

assign \reconfig_writedata[3]~input_o  = reconfig_writedata[3];

assign \reconfig_writedata[4]~input_o  = reconfig_writedata[4];

assign \reconfig_writedata[5]~input_o  = reconfig_writedata[5];

assign \reconfig_writedata[6]~input_o  = reconfig_writedata[6];

assign \reconfig_writedata[7]~input_o  = reconfig_writedata[7];

assign \rx_seriallpbken[0]~input_o  = rx_seriallpbken[0];

assign \tx_digitalreset[0]~input_o  = tx_digitalreset[0];

assign \tx_coreclkin[0]~input_o  = tx_coreclkin[0];

assign \tx_parallel_data[0]~input_o  = tx_parallel_data[0];

assign \tx_parallel_data[1]~input_o  = tx_parallel_data[1];

assign \tx_parallel_data[2]~input_o  = tx_parallel_data[2];

assign \tx_parallel_data[3]~input_o  = tx_parallel_data[3];

assign \tx_parallel_data[4]~input_o  = tx_parallel_data[4];

assign \tx_parallel_data[5]~input_o  = tx_parallel_data[5];

assign \tx_parallel_data[6]~input_o  = tx_parallel_data[6];

assign \tx_parallel_data[7]~input_o  = tx_parallel_data[7];

assign \tx_datak~input_o  = tx_datak;

assign \unused_tx_parallel_data[0]~input_o  = unused_tx_parallel_data[0];

assign \unused_tx_parallel_data[1]~input_o  = unused_tx_parallel_data[1];

assign \unused_tx_parallel_data[2]~input_o  = unused_tx_parallel_data[2];

assign \unused_tx_parallel_data[3]~input_o  = unused_tx_parallel_data[3];

assign \unused_tx_parallel_data[4]~input_o  = unused_tx_parallel_data[4];

assign \unused_tx_parallel_data[5]~input_o  = unused_tx_parallel_data[5];

assign \unused_tx_parallel_data[6]~input_o  = unused_tx_parallel_data[6];

assign \unused_tx_parallel_data[7]~input_o  = unused_tx_parallel_data[7];

assign \unused_tx_parallel_data[8]~input_o  = unused_tx_parallel_data[8];

assign \unused_tx_parallel_data[9]~input_o  = unused_tx_parallel_data[9];

assign \unused_tx_parallel_data[10]~input_o  = unused_tx_parallel_data[10];

assign \unused_tx_parallel_data[11]~input_o  = unused_tx_parallel_data[11];

assign \unused_tx_parallel_data[12]~input_o  = unused_tx_parallel_data[12];

assign \unused_tx_parallel_data[13]~input_o  = unused_tx_parallel_data[13];

assign \unused_tx_parallel_data[14]~input_o  = unused_tx_parallel_data[14];

assign \unused_tx_parallel_data[15]~input_o  = unused_tx_parallel_data[15];

assign \unused_tx_parallel_data[16]~input_o  = unused_tx_parallel_data[16];

assign \unused_tx_parallel_data[17]~input_o  = unused_tx_parallel_data[17];

assign \unused_tx_parallel_data[18]~input_o  = unused_tx_parallel_data[18];

assign \unused_tx_parallel_data[19]~input_o  = unused_tx_parallel_data[19];

assign \unused_tx_parallel_data[20]~input_o  = unused_tx_parallel_data[20];

assign \unused_tx_parallel_data[21]~input_o  = unused_tx_parallel_data[21];

assign \unused_tx_parallel_data[22]~input_o  = unused_tx_parallel_data[22];

assign \unused_tx_parallel_data[23]~input_o  = unused_tx_parallel_data[23];

assign \unused_tx_parallel_data[24]~input_o  = unused_tx_parallel_data[24];

assign \unused_tx_parallel_data[25]~input_o  = unused_tx_parallel_data[25];

assign \unused_tx_parallel_data[26]~input_o  = unused_tx_parallel_data[26];

assign \unused_tx_parallel_data[27]~input_o  = unused_tx_parallel_data[27];

assign \unused_tx_parallel_data[28]~input_o  = unused_tx_parallel_data[28];

assign \unused_tx_parallel_data[29]~input_o  = unused_tx_parallel_data[29];

assign \unused_tx_parallel_data[30]~input_o  = unused_tx_parallel_data[30];

assign \unused_tx_parallel_data[31]~input_o  = unused_tx_parallel_data[31];

assign \unused_tx_parallel_data[32]~input_o  = unused_tx_parallel_data[32];

assign \unused_tx_parallel_data[33]~input_o  = unused_tx_parallel_data[33];

assign \unused_tx_parallel_data[34]~input_o  = unused_tx_parallel_data[34];

assign \unused_tx_parallel_data[35]~input_o  = unused_tx_parallel_data[35];

assign \unused_tx_parallel_data[36]~input_o  = unused_tx_parallel_data[36];

assign \unused_tx_parallel_data[37]~input_o  = unused_tx_parallel_data[37];

assign \unused_tx_parallel_data[38]~input_o  = unused_tx_parallel_data[38];

assign \unused_tx_parallel_data[39]~input_o  = unused_tx_parallel_data[39];

assign \unused_tx_parallel_data[40]~input_o  = unused_tx_parallel_data[40];

assign \unused_tx_parallel_data[41]~input_o  = unused_tx_parallel_data[41];

assign \unused_tx_parallel_data[42]~input_o  = unused_tx_parallel_data[42];

assign \unused_tx_parallel_data[43]~input_o  = unused_tx_parallel_data[43];

assign \unused_tx_parallel_data[44]~input_o  = unused_tx_parallel_data[44];

assign \unused_tx_parallel_data[45]~input_o  = unused_tx_parallel_data[45];

assign \unused_tx_parallel_data[46]~input_o  = unused_tx_parallel_data[46];

assign \unused_tx_parallel_data[47]~input_o  = unused_tx_parallel_data[47];

assign \unused_tx_parallel_data[48]~input_o  = unused_tx_parallel_data[48];

assign \unused_tx_parallel_data[49]~input_o  = unused_tx_parallel_data[49];

assign \unused_tx_parallel_data[50]~input_o  = unused_tx_parallel_data[50];

assign \unused_tx_parallel_data[51]~input_o  = unused_tx_parallel_data[51];

assign \unused_tx_parallel_data[52]~input_o  = unused_tx_parallel_data[52];

assign \unused_tx_parallel_data[53]~input_o  = unused_tx_parallel_data[53];

assign \unused_tx_parallel_data[54]~input_o  = unused_tx_parallel_data[54];

assign \unused_tx_parallel_data[55]~input_o  = unused_tx_parallel_data[55];

assign \unused_tx_parallel_data[56]~input_o  = unused_tx_parallel_data[56];

assign \unused_tx_parallel_data[57]~input_o  = unused_tx_parallel_data[57];

assign \unused_tx_parallel_data[58]~input_o  = unused_tx_parallel_data[58];

assign \unused_tx_parallel_data[59]~input_o  = unused_tx_parallel_data[59];

assign \unused_tx_parallel_data[60]~input_o  = unused_tx_parallel_data[60];

assign \unused_tx_parallel_data[61]~input_o  = unused_tx_parallel_data[61];

assign \unused_tx_parallel_data[62]~input_o  = unused_tx_parallel_data[62];

assign \unused_tx_parallel_data[63]~input_o  = unused_tx_parallel_data[63];

assign \unused_tx_parallel_data[64]~input_o  = unused_tx_parallel_data[64];

assign \unused_tx_parallel_data[65]~input_o  = unused_tx_parallel_data[65];

assign \unused_tx_parallel_data[66]~input_o  = unused_tx_parallel_data[66];

assign \unused_tx_parallel_data[67]~input_o  = unused_tx_parallel_data[67];

assign \unused_tx_parallel_data[68]~input_o  = unused_tx_parallel_data[68];

assign \unused_tx_parallel_data[69]~input_o  = unused_tx_parallel_data[69];

assign \unused_tx_parallel_data[70]~input_o  = unused_tx_parallel_data[70];

assign \unused_tx_parallel_data[71]~input_o  = unused_tx_parallel_data[71];

assign \unused_tx_parallel_data[72]~input_o  = unused_tx_parallel_data[72];

assign \unused_tx_parallel_data[73]~input_o  = unused_tx_parallel_data[73];

assign \unused_tx_parallel_data[74]~input_o  = unused_tx_parallel_data[74];

assign \unused_tx_parallel_data[75]~input_o  = unused_tx_parallel_data[75];

assign \unused_tx_parallel_data[76]~input_o  = unused_tx_parallel_data[76];

assign \unused_tx_parallel_data[77]~input_o  = unused_tx_parallel_data[77];

assign \unused_tx_parallel_data[78]~input_o  = unused_tx_parallel_data[78];

assign \unused_tx_parallel_data[79]~input_o  = unused_tx_parallel_data[79];

assign \unused_tx_parallel_data[80]~input_o  = unused_tx_parallel_data[80];

assign \unused_tx_parallel_data[81]~input_o  = unused_tx_parallel_data[81];

assign \unused_tx_parallel_data[82]~input_o  = unused_tx_parallel_data[82];

assign \unused_tx_parallel_data[83]~input_o  = unused_tx_parallel_data[83];

assign \unused_tx_parallel_data[84]~input_o  = unused_tx_parallel_data[84];

assign \unused_tx_parallel_data[85]~input_o  = unused_tx_parallel_data[85];

assign \unused_tx_parallel_data[86]~input_o  = unused_tx_parallel_data[86];

assign \unused_tx_parallel_data[87]~input_o  = unused_tx_parallel_data[87];

assign \unused_tx_parallel_data[88]~input_o  = unused_tx_parallel_data[88];

assign \unused_tx_parallel_data[89]~input_o  = unused_tx_parallel_data[89];

assign \unused_tx_parallel_data[90]~input_o  = unused_tx_parallel_data[90];

assign \unused_tx_parallel_data[91]~input_o  = unused_tx_parallel_data[91];

assign \unused_tx_parallel_data[92]~input_o  = unused_tx_parallel_data[92];

assign \unused_tx_parallel_data[93]~input_o  = unused_tx_parallel_data[93];

assign \unused_tx_parallel_data[94]~input_o  = unused_tx_parallel_data[94];

assign \unused_tx_parallel_data[95]~input_o  = unused_tx_parallel_data[95];

assign \unused_tx_parallel_data[96]~input_o  = unused_tx_parallel_data[96];

assign \unused_tx_parallel_data[97]~input_o  = unused_tx_parallel_data[97];

assign \unused_tx_parallel_data[98]~input_o  = unused_tx_parallel_data[98];

assign \unused_tx_parallel_data[99]~input_o  = unused_tx_parallel_data[99];

assign \unused_tx_parallel_data[100]~input_o  = unused_tx_parallel_data[100];

assign \unused_tx_parallel_data[101]~input_o  = unused_tx_parallel_data[101];

assign \unused_tx_parallel_data[102]~input_o  = unused_tx_parallel_data[102];

assign \unused_tx_parallel_data[103]~input_o  = unused_tx_parallel_data[103];

assign \unused_tx_parallel_data[104]~input_o  = unused_tx_parallel_data[104];

assign \unused_tx_parallel_data[105]~input_o  = unused_tx_parallel_data[105];

assign \unused_tx_parallel_data[106]~input_o  = unused_tx_parallel_data[106];

assign \unused_tx_parallel_data[107]~input_o  = unused_tx_parallel_data[107];

assign \unused_tx_parallel_data[108]~input_o  = unused_tx_parallel_data[108];

assign \unused_tx_parallel_data[109]~input_o  = unused_tx_parallel_data[109];

assign \unused_tx_parallel_data[110]~input_o  = unused_tx_parallel_data[110];

assign \unused_tx_parallel_data[111]~input_o  = unused_tx_parallel_data[111];

assign \unused_tx_parallel_data[112]~input_o  = unused_tx_parallel_data[112];

assign \unused_tx_parallel_data[113]~input_o  = unused_tx_parallel_data[113];

assign \unused_tx_parallel_data[114]~input_o  = unused_tx_parallel_data[114];

assign \unused_tx_parallel_data[115]~input_o  = unused_tx_parallel_data[115];

assign \unused_tx_parallel_data[116]~input_o  = unused_tx_parallel_data[116];

assign \unused_tx_parallel_data[117]~input_o  = unused_tx_parallel_data[117];

assign \unused_tx_parallel_data[118]~input_o  = unused_tx_parallel_data[118];

assign \rx_serial_data[0]~input_o  = rx_serial_data[0];

assign \tx_serial_clk0[0]~input_o  = tx_serial_clk0[0];

assign \rx_cdr_refclk0~input_o  = rx_cdr_refclk0;

assign \reconfig_reset[0]~input_o  = reconfig_reset[0];

assign reconfig_readdata[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[0] ;

assign reconfig_readdata[1] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[1] ;

assign reconfig_readdata[2] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[2] ;

assign reconfig_readdata[3] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[3] ;

assign reconfig_readdata[4] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[4] ;

assign reconfig_readdata[5] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[5] ;

assign reconfig_readdata[6] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[6] ;

assign reconfig_readdata[7] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_readdata[7] ;

assign reconfig_readdata[8] = gnd;

assign reconfig_readdata[9] = gnd;

assign reconfig_readdata[10] = gnd;

assign reconfig_readdata[11] = gnd;

assign reconfig_readdata[12] = gnd;

assign reconfig_readdata[13] = gnd;

assign reconfig_readdata[14] = gnd;

assign reconfig_readdata[15] = gnd;

assign reconfig_readdata[16] = gnd;

assign reconfig_readdata[17] = gnd;

assign reconfig_readdata[18] = gnd;

assign reconfig_readdata[19] = gnd;

assign reconfig_readdata[20] = gnd;

assign reconfig_readdata[21] = gnd;

assign reconfig_readdata[22] = gnd;

assign reconfig_readdata[23] = gnd;

assign reconfig_readdata[24] = gnd;

assign reconfig_readdata[25] = gnd;

assign reconfig_readdata[26] = gnd;

assign reconfig_readdata[27] = gnd;

assign reconfig_readdata[28] = gnd;

assign reconfig_readdata[29] = gnd;

assign reconfig_readdata[30] = gnd;

assign reconfig_readdata[31] = gnd;

assign reconfig_waitrequest[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|avmm_waitrequest[0]~0_combout ;

assign rx_cal_busy[0] = ~ \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|pld_cal_done[0] ;

assign rx_clkout[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out ;

assign rx_datak = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[8] ;

assign rx_disperr = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[11] ;

assign rx_errdetect = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[9] ;

assign rx_is_lockedtodata[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock ;

assign rx_is_lockedtoref[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock ;

assign rx_parallel_data[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[0] ;

assign rx_parallel_data[1] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[1] ;

assign rx_parallel_data[2] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[2] ;

assign rx_parallel_data[3] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[3] ;

assign rx_parallel_data[4] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[4] ;

assign rx_parallel_data[5] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[5] ;

assign rx_parallel_data[6] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[6] ;

assign rx_parallel_data[7] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[7] ;

assign rx_patterndetect = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[12] ;

assign rx_runningdisp = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[15] ;

assign rx_std_bitslipboundarysel[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[0] ;

assign rx_std_bitslipboundarysel[1] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[1] ;

assign rx_std_bitslipboundarysel[2] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[2] ;

assign rx_std_bitslipboundarysel[3] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[3] ;

assign rx_std_bitslipboundarysel[4] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary[4] ;

assign rx_syncstatus = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[10] ;

assign tx_cal_busy[0] = ~ \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_xcvr_avmm|pld_cal_done[0] ;

assign tx_clkout[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_pld_pcs_tx_clk_out ;

assign tx_serial_data[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pma|w_pma_tx_buf_vop ;

assign unused_rx_parallel_data[0] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[13] ;

assign unused_rx_parallel_data[1] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[14] ;

assign unused_rx_parallel_data[2] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[16] ;

assign unused_rx_parallel_data[3] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[17] ;

assign unused_rx_parallel_data[4] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[18] ;

assign unused_rx_parallel_data[5] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[19] ;

assign unused_rx_parallel_data[6] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[20] ;

assign unused_rx_parallel_data[7] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[21] ;

assign unused_rx_parallel_data[8] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[22] ;

assign unused_rx_parallel_data[9] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[23] ;

assign unused_rx_parallel_data[10] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[24] ;

assign unused_rx_parallel_data[11] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[25] ;

assign unused_rx_parallel_data[12] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[26] ;

assign unused_rx_parallel_data[13] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[27] ;

assign unused_rx_parallel_data[14] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[28] ;

assign unused_rx_parallel_data[15] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[29] ;

assign unused_rx_parallel_data[16] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[30] ;

assign unused_rx_parallel_data[17] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[31] ;

assign unused_rx_parallel_data[18] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[32] ;

assign unused_rx_parallel_data[19] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[33] ;

assign unused_rx_parallel_data[20] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[34] ;

assign unused_rx_parallel_data[21] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[35] ;

assign unused_rx_parallel_data[22] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[36] ;

assign unused_rx_parallel_data[23] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[37] ;

assign unused_rx_parallel_data[24] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[38] ;

assign unused_rx_parallel_data[25] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[39] ;

assign unused_rx_parallel_data[26] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[40] ;

assign unused_rx_parallel_data[27] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[41] ;

assign unused_rx_parallel_data[28] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[42] ;

assign unused_rx_parallel_data[29] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[43] ;

assign unused_rx_parallel_data[30] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[44] ;

assign unused_rx_parallel_data[31] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[45] ;

assign unused_rx_parallel_data[32] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[46] ;

assign unused_rx_parallel_data[33] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[47] ;

assign unused_rx_parallel_data[34] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[48] ;

assign unused_rx_parallel_data[35] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[49] ;

assign unused_rx_parallel_data[36] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[50] ;

assign unused_rx_parallel_data[37] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[51] ;

assign unused_rx_parallel_data[38] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[52] ;

assign unused_rx_parallel_data[39] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[53] ;

assign unused_rx_parallel_data[40] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[54] ;

assign unused_rx_parallel_data[41] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[55] ;

assign unused_rx_parallel_data[42] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[56] ;

assign unused_rx_parallel_data[43] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[57] ;

assign unused_rx_parallel_data[44] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[58] ;

assign unused_rx_parallel_data[45] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[59] ;

assign unused_rx_parallel_data[46] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[60] ;

assign unused_rx_parallel_data[47] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[61] ;

assign unused_rx_parallel_data[48] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[62] ;

assign unused_rx_parallel_data[49] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[63] ;

assign unused_rx_parallel_data[50] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[64] ;

assign unused_rx_parallel_data[51] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[65] ;

assign unused_rx_parallel_data[52] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[66] ;

assign unused_rx_parallel_data[53] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[67] ;

assign unused_rx_parallel_data[54] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[68] ;

assign unused_rx_parallel_data[55] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[69] ;

assign unused_rx_parallel_data[56] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[70] ;

assign unused_rx_parallel_data[57] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[71] ;

assign unused_rx_parallel_data[58] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[72] ;

assign unused_rx_parallel_data[59] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[73] ;

assign unused_rx_parallel_data[60] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[74] ;

assign unused_rx_parallel_data[61] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[75] ;

assign unused_rx_parallel_data[62] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[76] ;

assign unused_rx_parallel_data[63] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[77] ;

assign unused_rx_parallel_data[64] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[78] ;

assign unused_rx_parallel_data[65] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[79] ;

assign unused_rx_parallel_data[66] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[80] ;

assign unused_rx_parallel_data[67] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[81] ;

assign unused_rx_parallel_data[68] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[82] ;

assign unused_rx_parallel_data[69] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[83] ;

assign unused_rx_parallel_data[70] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[84] ;

assign unused_rx_parallel_data[71] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[85] ;

assign unused_rx_parallel_data[72] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[86] ;

assign unused_rx_parallel_data[73] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[87] ;

assign unused_rx_parallel_data[74] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[88] ;

assign unused_rx_parallel_data[75] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[89] ;

assign unused_rx_parallel_data[76] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[90] ;

assign unused_rx_parallel_data[77] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[91] ;

assign unused_rx_parallel_data[78] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[92] ;

assign unused_rx_parallel_data[79] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[93] ;

assign unused_rx_parallel_data[80] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[94] ;

assign unused_rx_parallel_data[81] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[95] ;

assign unused_rx_parallel_data[82] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[96] ;

assign unused_rx_parallel_data[83] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[97] ;

assign unused_rx_parallel_data[84] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[98] ;

assign unused_rx_parallel_data[85] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[99] ;

assign unused_rx_parallel_data[86] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[100] ;

assign unused_rx_parallel_data[87] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[101] ;

assign unused_rx_parallel_data[88] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[102] ;

assign unused_rx_parallel_data[89] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[103] ;

assign unused_rx_parallel_data[90] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[104] ;

assign unused_rx_parallel_data[91] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[105] ;

assign unused_rx_parallel_data[92] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[106] ;

assign unused_rx_parallel_data[93] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[107] ;

assign unused_rx_parallel_data[94] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[108] ;

assign unused_rx_parallel_data[95] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[109] ;

assign unused_rx_parallel_data[96] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[110] ;

assign unused_rx_parallel_data[97] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[111] ;

assign unused_rx_parallel_data[98] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[112] ;

assign unused_rx_parallel_data[99] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[113] ;

assign unused_rx_parallel_data[100] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[114] ;

assign unused_rx_parallel_data[101] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[115] ;

assign unused_rx_parallel_data[102] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[116] ;

assign unused_rx_parallel_data[103] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[117] ;

assign unused_rx_parallel_data[104] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[118] ;

assign unused_rx_parallel_data[105] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[119] ;

assign unused_rx_parallel_data[106] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[120] ;

assign unused_rx_parallel_data[107] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[121] ;

assign unused_rx_parallel_data[108] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[122] ;

assign unused_rx_parallel_data[109] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[123] ;

assign unused_rx_parallel_data[110] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[124] ;

assign unused_rx_parallel_data[111] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[125] ;

assign unused_rx_parallel_data[112] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[126] ;

assign unused_rx_parallel_data[113] = \xcvr_native_a10_0|g_xcvr_native_insts[0].twentynm_xcvr_native_inst|twentynm_xcvr_native_inst|inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_pld_rx_data[127] ;

twentynm_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

assign \reconfig_address[9]~input_o  = reconfig_address[9];

assign \reconfig_writedata[8]~input_o  = reconfig_writedata[8];

assign \reconfig_writedata[9]~input_o  = reconfig_writedata[9];

assign \reconfig_writedata[10]~input_o  = reconfig_writedata[10];

assign \reconfig_writedata[11]~input_o  = reconfig_writedata[11];

assign \reconfig_writedata[12]~input_o  = reconfig_writedata[12];

assign \reconfig_writedata[13]~input_o  = reconfig_writedata[13];

assign \reconfig_writedata[14]~input_o  = reconfig_writedata[14];

assign \reconfig_writedata[15]~input_o  = reconfig_writedata[15];

assign \reconfig_writedata[16]~input_o  = reconfig_writedata[16];

assign \reconfig_writedata[17]~input_o  = reconfig_writedata[17];

assign \reconfig_writedata[18]~input_o  = reconfig_writedata[18];

assign \reconfig_writedata[19]~input_o  = reconfig_writedata[19];

assign \reconfig_writedata[20]~input_o  = reconfig_writedata[20];

assign \reconfig_writedata[21]~input_o  = reconfig_writedata[21];

assign \reconfig_writedata[22]~input_o  = reconfig_writedata[22];

assign \reconfig_writedata[23]~input_o  = reconfig_writedata[23];

assign \reconfig_writedata[24]~input_o  = reconfig_writedata[24];

assign \reconfig_writedata[25]~input_o  = reconfig_writedata[25];

assign \reconfig_writedata[26]~input_o  = reconfig_writedata[26];

assign \reconfig_writedata[27]~input_o  = reconfig_writedata[27];

assign \reconfig_writedata[28]~input_o  = reconfig_writedata[28];

assign \reconfig_writedata[29]~input_o  = reconfig_writedata[29];

assign \reconfig_writedata[30]~input_o  = reconfig_writedata[30];

assign \reconfig_writedata[31]~input_o  = reconfig_writedata[31];

endmodule

module wr_arria10_e3p1_det_phy_wr_arria10_e3p1_det_phy_altera_xcvr_native_a10_181_iwfuxyq (
	w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_0,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_1,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_2,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_3,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_5,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_6,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_7,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_8,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_9,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_10,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_11,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_12,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_13,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_14,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_15,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_16,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_17,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_18,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_19,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_20,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_21,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_22,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_23,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_24,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_25,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_26,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_27,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_28,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_29,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_30,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_31,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_32,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_33,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_34,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_35,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_36,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_37,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_38,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_39,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_40,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_41,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_42,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_43,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_44,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_45,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_46,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_47,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_48,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_49,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_50,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_51,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_52,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_53,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_54,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_55,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_56,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_57,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_58,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_59,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_60,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_61,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_62,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_63,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_64,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_65,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_66,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_67,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_68,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_69,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_70,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_71,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_72,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_73,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_74,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_75,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_76,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_77,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_78,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_79,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_80,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_81,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_82,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_83,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_84,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_85,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_86,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_87,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_88,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_89,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_90,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_91,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_92,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_93,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_94,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_95,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_96,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_97,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_98,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_99,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_100,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_101,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_102,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_103,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_104,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_105,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_106,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_107,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_108,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_109,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_110,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_111,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_112,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_113,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_114,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_115,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_116,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_117,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_118,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_119,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_120,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_121,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_122,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_123,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_124,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_125,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_126,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_127,
	pld_cal_done_0,
	avmm_readdata_0,
	avmm_readdata_1,
	avmm_readdata_2,
	avmm_readdata_3,
	avmm_readdata_4,
	avmm_readdata_5,
	avmm_readdata_6,
	avmm_readdata_7,
	w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock,
	w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock,
	tx_clkout,
	tx_serial_data,
	avmm_waitrequest_0,
	reset_out_stage_0,
	reset_out_stage_1,
	reconfig_read_0,
	rx_digitalreset_0,
	rx_std_wa_patternalign_0,
	rx_coreclkin_0,
	reconfig_clk_0,
	reconfig_write_0,
	reconfig_address_0,
	reconfig_address_1,
	reconfig_address_2,
	reconfig_address_3,
	reconfig_address_4,
	reconfig_address_5,
	reconfig_address_6,
	reconfig_address_7,
	reconfig_address_8,
	reconfig_writedata_0,
	reconfig_writedata_1,
	reconfig_writedata_2,
	reconfig_writedata_3,
	reconfig_writedata_4,
	reconfig_writedata_5,
	reconfig_writedata_6,
	reconfig_writedata_7,
	rx_seriallpbken_0,
	tx_digitalreset_0,
	tx_coreclkin_0,
	tx_parallel_data_0,
	tx_parallel_data_1,
	tx_parallel_data_2,
	tx_parallel_data_3,
	tx_parallel_data_4,
	tx_parallel_data_5,
	tx_parallel_data_6,
	tx_parallel_data_7,
	tx_datak,
	unused_tx_parallel_data_0,
	unused_tx_parallel_data_1,
	unused_tx_parallel_data_2,
	unused_tx_parallel_data_3,
	unused_tx_parallel_data_4,
	unused_tx_parallel_data_5,
	unused_tx_parallel_data_6,
	unused_tx_parallel_data_7,
	unused_tx_parallel_data_8,
	unused_tx_parallel_data_9,
	unused_tx_parallel_data_10,
	unused_tx_parallel_data_11,
	unused_tx_parallel_data_12,
	unused_tx_parallel_data_13,
	unused_tx_parallel_data_14,
	unused_tx_parallel_data_15,
	unused_tx_parallel_data_16,
	unused_tx_parallel_data_17,
	unused_tx_parallel_data_18,
	unused_tx_parallel_data_19,
	unused_tx_parallel_data_20,
	unused_tx_parallel_data_21,
	unused_tx_parallel_data_22,
	unused_tx_parallel_data_23,
	unused_tx_parallel_data_24,
	unused_tx_parallel_data_25,
	unused_tx_parallel_data_26,
	unused_tx_parallel_data_27,
	unused_tx_parallel_data_28,
	unused_tx_parallel_data_29,
	unused_tx_parallel_data_30,
	unused_tx_parallel_data_31,
	unused_tx_parallel_data_32,
	unused_tx_parallel_data_33,
	unused_tx_parallel_data_34,
	unused_tx_parallel_data_35,
	unused_tx_parallel_data_36,
	unused_tx_parallel_data_37,
	unused_tx_parallel_data_38,
	unused_tx_parallel_data_39,
	unused_tx_parallel_data_40,
	unused_tx_parallel_data_41,
	unused_tx_parallel_data_42,
	unused_tx_parallel_data_43,
	unused_tx_parallel_data_44,
	unused_tx_parallel_data_45,
	unused_tx_parallel_data_46,
	unused_tx_parallel_data_47,
	unused_tx_parallel_data_48,
	unused_tx_parallel_data_49,
	unused_tx_parallel_data_50,
	unused_tx_parallel_data_51,
	unused_tx_parallel_data_52,
	unused_tx_parallel_data_53,
	unused_tx_parallel_data_54,
	unused_tx_parallel_data_55,
	unused_tx_parallel_data_56,
	unused_tx_parallel_data_57,
	unused_tx_parallel_data_58,
	unused_tx_parallel_data_59,
	unused_tx_parallel_data_60,
	unused_tx_parallel_data_61,
	unused_tx_parallel_data_62,
	unused_tx_parallel_data_63,
	unused_tx_parallel_data_64,
	unused_tx_parallel_data_65,
	unused_tx_parallel_data_66,
	unused_tx_parallel_data_67,
	unused_tx_parallel_data_68,
	unused_tx_parallel_data_69,
	unused_tx_parallel_data_70,
	unused_tx_parallel_data_71,
	unused_tx_parallel_data_72,
	unused_tx_parallel_data_73,
	unused_tx_parallel_data_74,
	unused_tx_parallel_data_75,
	unused_tx_parallel_data_76,
	unused_tx_parallel_data_77,
	unused_tx_parallel_data_78,
	unused_tx_parallel_data_79,
	unused_tx_parallel_data_80,
	unused_tx_parallel_data_81,
	unused_tx_parallel_data_82,
	unused_tx_parallel_data_83,
	unused_tx_parallel_data_84,
	unused_tx_parallel_data_85,
	unused_tx_parallel_data_86,
	unused_tx_parallel_data_87,
	unused_tx_parallel_data_88,
	unused_tx_parallel_data_89,
	unused_tx_parallel_data_90,
	unused_tx_parallel_data_91,
	unused_tx_parallel_data_92,
	unused_tx_parallel_data_93,
	unused_tx_parallel_data_94,
	unused_tx_parallel_data_95,
	unused_tx_parallel_data_96,
	unused_tx_parallel_data_97,
	unused_tx_parallel_data_98,
	unused_tx_parallel_data_99,
	unused_tx_parallel_data_100,
	unused_tx_parallel_data_101,
	unused_tx_parallel_data_102,
	unused_tx_parallel_data_103,
	unused_tx_parallel_data_104,
	unused_tx_parallel_data_105,
	unused_tx_parallel_data_106,
	unused_tx_parallel_data_107,
	unused_tx_parallel_data_108,
	unused_tx_parallel_data_109,
	unused_tx_parallel_data_110,
	unused_tx_parallel_data_111,
	unused_tx_parallel_data_112,
	unused_tx_parallel_data_113,
	unused_tx_parallel_data_114,
	unused_tx_parallel_data_115,
	unused_tx_parallel_data_116,
	unused_tx_parallel_data_117,
	unused_tx_parallel_data_118,
	rx_serial_data_0,
	tx_serial_clk0_0,
	rx_cdr_refclk0,
	reconfig_reset_0)/* synthesis synthesis_greybox=1 */;
output 	w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_0;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_1;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_2;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_3;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_5;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_6;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_7;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_8;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_9;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_10;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_11;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_12;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_13;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_14;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_15;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_16;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_17;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_18;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_19;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_20;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_21;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_22;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_23;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_24;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_25;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_26;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_27;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_28;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_29;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_30;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_31;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_32;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_33;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_34;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_35;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_36;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_37;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_38;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_39;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_40;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_41;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_42;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_43;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_44;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_45;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_46;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_47;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_48;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_49;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_50;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_51;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_52;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_53;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_54;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_55;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_56;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_57;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_58;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_59;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_60;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_61;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_62;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_63;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_64;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_65;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_66;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_67;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_68;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_69;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_70;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_71;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_72;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_73;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_74;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_75;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_76;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_77;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_78;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_79;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_80;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_81;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_82;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_83;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_84;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_85;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_86;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_87;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_88;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_89;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_90;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_91;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_92;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_93;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_94;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_95;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_96;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_97;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_98;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_99;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_100;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_101;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_102;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_103;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_104;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_105;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_106;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_107;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_108;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_109;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_110;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_111;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_112;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_113;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_114;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_115;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_116;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_117;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_118;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_119;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_120;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_121;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_122;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_123;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_124;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_125;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_126;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_127;
output 	pld_cal_done_0;
output 	avmm_readdata_0;
output 	avmm_readdata_1;
output 	avmm_readdata_2;
output 	avmm_readdata_3;
output 	avmm_readdata_4;
output 	avmm_readdata_5;
output 	avmm_readdata_6;
output 	avmm_readdata_7;
output 	w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock;
output 	w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock;
output 	[0:0] tx_clkout;
output 	[0:0] tx_serial_data;
output 	avmm_waitrequest_0;
input 	reset_out_stage_0;
input 	reset_out_stage_1;
input 	reconfig_read_0;
input 	rx_digitalreset_0;
input 	rx_std_wa_patternalign_0;
input 	rx_coreclkin_0;
input 	reconfig_clk_0;
input 	reconfig_write_0;
input 	reconfig_address_0;
input 	reconfig_address_1;
input 	reconfig_address_2;
input 	reconfig_address_3;
input 	reconfig_address_4;
input 	reconfig_address_5;
input 	reconfig_address_6;
input 	reconfig_address_7;
input 	reconfig_address_8;
input 	reconfig_writedata_0;
input 	reconfig_writedata_1;
input 	reconfig_writedata_2;
input 	reconfig_writedata_3;
input 	reconfig_writedata_4;
input 	reconfig_writedata_5;
input 	reconfig_writedata_6;
input 	reconfig_writedata_7;
input 	rx_seriallpbken_0;
input 	tx_digitalreset_0;
input 	tx_coreclkin_0;
input 	tx_parallel_data_0;
input 	tx_parallel_data_1;
input 	tx_parallel_data_2;
input 	tx_parallel_data_3;
input 	tx_parallel_data_4;
input 	tx_parallel_data_5;
input 	tx_parallel_data_6;
input 	tx_parallel_data_7;
input 	tx_datak;
input 	unused_tx_parallel_data_0;
input 	unused_tx_parallel_data_1;
input 	unused_tx_parallel_data_2;
input 	unused_tx_parallel_data_3;
input 	unused_tx_parallel_data_4;
input 	unused_tx_parallel_data_5;
input 	unused_tx_parallel_data_6;
input 	unused_tx_parallel_data_7;
input 	unused_tx_parallel_data_8;
input 	unused_tx_parallel_data_9;
input 	unused_tx_parallel_data_10;
input 	unused_tx_parallel_data_11;
input 	unused_tx_parallel_data_12;
input 	unused_tx_parallel_data_13;
input 	unused_tx_parallel_data_14;
input 	unused_tx_parallel_data_15;
input 	unused_tx_parallel_data_16;
input 	unused_tx_parallel_data_17;
input 	unused_tx_parallel_data_18;
input 	unused_tx_parallel_data_19;
input 	unused_tx_parallel_data_20;
input 	unused_tx_parallel_data_21;
input 	unused_tx_parallel_data_22;
input 	unused_tx_parallel_data_23;
input 	unused_tx_parallel_data_24;
input 	unused_tx_parallel_data_25;
input 	unused_tx_parallel_data_26;
input 	unused_tx_parallel_data_27;
input 	unused_tx_parallel_data_28;
input 	unused_tx_parallel_data_29;
input 	unused_tx_parallel_data_30;
input 	unused_tx_parallel_data_31;
input 	unused_tx_parallel_data_32;
input 	unused_tx_parallel_data_33;
input 	unused_tx_parallel_data_34;
input 	unused_tx_parallel_data_35;
input 	unused_tx_parallel_data_36;
input 	unused_tx_parallel_data_37;
input 	unused_tx_parallel_data_38;
input 	unused_tx_parallel_data_39;
input 	unused_tx_parallel_data_40;
input 	unused_tx_parallel_data_41;
input 	unused_tx_parallel_data_42;
input 	unused_tx_parallel_data_43;
input 	unused_tx_parallel_data_44;
input 	unused_tx_parallel_data_45;
input 	unused_tx_parallel_data_46;
input 	unused_tx_parallel_data_47;
input 	unused_tx_parallel_data_48;
input 	unused_tx_parallel_data_49;
input 	unused_tx_parallel_data_50;
input 	unused_tx_parallel_data_51;
input 	unused_tx_parallel_data_52;
input 	unused_tx_parallel_data_53;
input 	unused_tx_parallel_data_54;
input 	unused_tx_parallel_data_55;
input 	unused_tx_parallel_data_56;
input 	unused_tx_parallel_data_57;
input 	unused_tx_parallel_data_58;
input 	unused_tx_parallel_data_59;
input 	unused_tx_parallel_data_60;
input 	unused_tx_parallel_data_61;
input 	unused_tx_parallel_data_62;
input 	unused_tx_parallel_data_63;
input 	unused_tx_parallel_data_64;
input 	unused_tx_parallel_data_65;
input 	unused_tx_parallel_data_66;
input 	unused_tx_parallel_data_67;
input 	unused_tx_parallel_data_68;
input 	unused_tx_parallel_data_69;
input 	unused_tx_parallel_data_70;
input 	unused_tx_parallel_data_71;
input 	unused_tx_parallel_data_72;
input 	unused_tx_parallel_data_73;
input 	unused_tx_parallel_data_74;
input 	unused_tx_parallel_data_75;
input 	unused_tx_parallel_data_76;
input 	unused_tx_parallel_data_77;
input 	unused_tx_parallel_data_78;
input 	unused_tx_parallel_data_79;
input 	unused_tx_parallel_data_80;
input 	unused_tx_parallel_data_81;
input 	unused_tx_parallel_data_82;
input 	unused_tx_parallel_data_83;
input 	unused_tx_parallel_data_84;
input 	unused_tx_parallel_data_85;
input 	unused_tx_parallel_data_86;
input 	unused_tx_parallel_data_87;
input 	unused_tx_parallel_data_88;
input 	unused_tx_parallel_data_89;
input 	unused_tx_parallel_data_90;
input 	unused_tx_parallel_data_91;
input 	unused_tx_parallel_data_92;
input 	unused_tx_parallel_data_93;
input 	unused_tx_parallel_data_94;
input 	unused_tx_parallel_data_95;
input 	unused_tx_parallel_data_96;
input 	unused_tx_parallel_data_97;
input 	unused_tx_parallel_data_98;
input 	unused_tx_parallel_data_99;
input 	unused_tx_parallel_data_100;
input 	unused_tx_parallel_data_101;
input 	unused_tx_parallel_data_102;
input 	unused_tx_parallel_data_103;
input 	unused_tx_parallel_data_104;
input 	unused_tx_parallel_data_105;
input 	unused_tx_parallel_data_106;
input 	unused_tx_parallel_data_107;
input 	unused_tx_parallel_data_108;
input 	unused_tx_parallel_data_109;
input 	unused_tx_parallel_data_110;
input 	unused_tx_parallel_data_111;
input 	unused_tx_parallel_data_112;
input 	unused_tx_parallel_data_113;
input 	unused_tx_parallel_data_114;
input 	unused_tx_parallel_data_115;
input 	unused_tx_parallel_data_116;
input 	unused_tx_parallel_data_117;
input 	unused_tx_parallel_data_118;
input 	rx_serial_data_0;
input 	tx_serial_clk0_0;
input 	rx_cdr_refclk0;
input 	reconfig_reset_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



wr_arria10_e3p1_det_phy_twentynm_xcvr_native \g_xcvr_native_insts[0].twentynm_xcvr_native_inst (
	.out_pld_pcs_rx_clk_out(w_hssi_rx_pld_pcs_interface_pld_pcs_rx_clk_out),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_0(w_hssi_rx_pld_pcs_interface_pld_rx_data_0),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_1(w_hssi_rx_pld_pcs_interface_pld_rx_data_1),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_2(w_hssi_rx_pld_pcs_interface_pld_rx_data_2),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_3(w_hssi_rx_pld_pcs_interface_pld_rx_data_3),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_4(w_hssi_rx_pld_pcs_interface_pld_rx_data_4),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_5(w_hssi_rx_pld_pcs_interface_pld_rx_data_5),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_6(w_hssi_rx_pld_pcs_interface_pld_rx_data_6),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_7(w_hssi_rx_pld_pcs_interface_pld_rx_data_7),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_8(w_hssi_rx_pld_pcs_interface_pld_rx_data_8),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_9(w_hssi_rx_pld_pcs_interface_pld_rx_data_9),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_10(w_hssi_rx_pld_pcs_interface_pld_rx_data_10),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_11(w_hssi_rx_pld_pcs_interface_pld_rx_data_11),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_12(w_hssi_rx_pld_pcs_interface_pld_rx_data_12),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_13(w_hssi_rx_pld_pcs_interface_pld_rx_data_13),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_14(w_hssi_rx_pld_pcs_interface_pld_rx_data_14),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_15(w_hssi_rx_pld_pcs_interface_pld_rx_data_15),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_16(w_hssi_rx_pld_pcs_interface_pld_rx_data_16),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_17(w_hssi_rx_pld_pcs_interface_pld_rx_data_17),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_18(w_hssi_rx_pld_pcs_interface_pld_rx_data_18),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_19(w_hssi_rx_pld_pcs_interface_pld_rx_data_19),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_20(w_hssi_rx_pld_pcs_interface_pld_rx_data_20),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_21(w_hssi_rx_pld_pcs_interface_pld_rx_data_21),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_22(w_hssi_rx_pld_pcs_interface_pld_rx_data_22),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_23(w_hssi_rx_pld_pcs_interface_pld_rx_data_23),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_24(w_hssi_rx_pld_pcs_interface_pld_rx_data_24),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_25(w_hssi_rx_pld_pcs_interface_pld_rx_data_25),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_26(w_hssi_rx_pld_pcs_interface_pld_rx_data_26),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_27(w_hssi_rx_pld_pcs_interface_pld_rx_data_27),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_28(w_hssi_rx_pld_pcs_interface_pld_rx_data_28),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_29(w_hssi_rx_pld_pcs_interface_pld_rx_data_29),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_30(w_hssi_rx_pld_pcs_interface_pld_rx_data_30),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_31(w_hssi_rx_pld_pcs_interface_pld_rx_data_31),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_32(w_hssi_rx_pld_pcs_interface_pld_rx_data_32),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_33(w_hssi_rx_pld_pcs_interface_pld_rx_data_33),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_34(w_hssi_rx_pld_pcs_interface_pld_rx_data_34),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_35(w_hssi_rx_pld_pcs_interface_pld_rx_data_35),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_36(w_hssi_rx_pld_pcs_interface_pld_rx_data_36),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_37(w_hssi_rx_pld_pcs_interface_pld_rx_data_37),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_38(w_hssi_rx_pld_pcs_interface_pld_rx_data_38),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_39(w_hssi_rx_pld_pcs_interface_pld_rx_data_39),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_40(w_hssi_rx_pld_pcs_interface_pld_rx_data_40),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_41(w_hssi_rx_pld_pcs_interface_pld_rx_data_41),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_42(w_hssi_rx_pld_pcs_interface_pld_rx_data_42),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_43(w_hssi_rx_pld_pcs_interface_pld_rx_data_43),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_44(w_hssi_rx_pld_pcs_interface_pld_rx_data_44),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_45(w_hssi_rx_pld_pcs_interface_pld_rx_data_45),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_46(w_hssi_rx_pld_pcs_interface_pld_rx_data_46),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_47(w_hssi_rx_pld_pcs_interface_pld_rx_data_47),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_48(w_hssi_rx_pld_pcs_interface_pld_rx_data_48),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_49(w_hssi_rx_pld_pcs_interface_pld_rx_data_49),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_50(w_hssi_rx_pld_pcs_interface_pld_rx_data_50),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_51(w_hssi_rx_pld_pcs_interface_pld_rx_data_51),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_52(w_hssi_rx_pld_pcs_interface_pld_rx_data_52),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_53(w_hssi_rx_pld_pcs_interface_pld_rx_data_53),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_54(w_hssi_rx_pld_pcs_interface_pld_rx_data_54),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_55(w_hssi_rx_pld_pcs_interface_pld_rx_data_55),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_56(w_hssi_rx_pld_pcs_interface_pld_rx_data_56),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_57(w_hssi_rx_pld_pcs_interface_pld_rx_data_57),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_58(w_hssi_rx_pld_pcs_interface_pld_rx_data_58),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_59(w_hssi_rx_pld_pcs_interface_pld_rx_data_59),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_60(w_hssi_rx_pld_pcs_interface_pld_rx_data_60),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_61(w_hssi_rx_pld_pcs_interface_pld_rx_data_61),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_62(w_hssi_rx_pld_pcs_interface_pld_rx_data_62),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_63(w_hssi_rx_pld_pcs_interface_pld_rx_data_63),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_64(w_hssi_rx_pld_pcs_interface_pld_rx_data_64),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_65(w_hssi_rx_pld_pcs_interface_pld_rx_data_65),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_66(w_hssi_rx_pld_pcs_interface_pld_rx_data_66),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_67(w_hssi_rx_pld_pcs_interface_pld_rx_data_67),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_68(w_hssi_rx_pld_pcs_interface_pld_rx_data_68),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_69(w_hssi_rx_pld_pcs_interface_pld_rx_data_69),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_70(w_hssi_rx_pld_pcs_interface_pld_rx_data_70),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_71(w_hssi_rx_pld_pcs_interface_pld_rx_data_71),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_72(w_hssi_rx_pld_pcs_interface_pld_rx_data_72),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_73(w_hssi_rx_pld_pcs_interface_pld_rx_data_73),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_74(w_hssi_rx_pld_pcs_interface_pld_rx_data_74),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_75(w_hssi_rx_pld_pcs_interface_pld_rx_data_75),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_76(w_hssi_rx_pld_pcs_interface_pld_rx_data_76),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_77(w_hssi_rx_pld_pcs_interface_pld_rx_data_77),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_78(w_hssi_rx_pld_pcs_interface_pld_rx_data_78),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_79(w_hssi_rx_pld_pcs_interface_pld_rx_data_79),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_80(w_hssi_rx_pld_pcs_interface_pld_rx_data_80),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_81(w_hssi_rx_pld_pcs_interface_pld_rx_data_81),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_82(w_hssi_rx_pld_pcs_interface_pld_rx_data_82),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_83(w_hssi_rx_pld_pcs_interface_pld_rx_data_83),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_84(w_hssi_rx_pld_pcs_interface_pld_rx_data_84),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_85(w_hssi_rx_pld_pcs_interface_pld_rx_data_85),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_86(w_hssi_rx_pld_pcs_interface_pld_rx_data_86),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_87(w_hssi_rx_pld_pcs_interface_pld_rx_data_87),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_88(w_hssi_rx_pld_pcs_interface_pld_rx_data_88),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_89(w_hssi_rx_pld_pcs_interface_pld_rx_data_89),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_90(w_hssi_rx_pld_pcs_interface_pld_rx_data_90),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_91(w_hssi_rx_pld_pcs_interface_pld_rx_data_91),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_92(w_hssi_rx_pld_pcs_interface_pld_rx_data_92),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_93(w_hssi_rx_pld_pcs_interface_pld_rx_data_93),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_94(w_hssi_rx_pld_pcs_interface_pld_rx_data_94),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_95(w_hssi_rx_pld_pcs_interface_pld_rx_data_95),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_96(w_hssi_rx_pld_pcs_interface_pld_rx_data_96),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_97(w_hssi_rx_pld_pcs_interface_pld_rx_data_97),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_98(w_hssi_rx_pld_pcs_interface_pld_rx_data_98),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_99(w_hssi_rx_pld_pcs_interface_pld_rx_data_99),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_100(w_hssi_rx_pld_pcs_interface_pld_rx_data_100),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_101(w_hssi_rx_pld_pcs_interface_pld_rx_data_101),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_102(w_hssi_rx_pld_pcs_interface_pld_rx_data_102),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_103(w_hssi_rx_pld_pcs_interface_pld_rx_data_103),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_104(w_hssi_rx_pld_pcs_interface_pld_rx_data_104),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_105(w_hssi_rx_pld_pcs_interface_pld_rx_data_105),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_106(w_hssi_rx_pld_pcs_interface_pld_rx_data_106),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_107(w_hssi_rx_pld_pcs_interface_pld_rx_data_107),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_108(w_hssi_rx_pld_pcs_interface_pld_rx_data_108),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_109(w_hssi_rx_pld_pcs_interface_pld_rx_data_109),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_110(w_hssi_rx_pld_pcs_interface_pld_rx_data_110),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_111(w_hssi_rx_pld_pcs_interface_pld_rx_data_111),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_112(w_hssi_rx_pld_pcs_interface_pld_rx_data_112),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_113(w_hssi_rx_pld_pcs_interface_pld_rx_data_113),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_114(w_hssi_rx_pld_pcs_interface_pld_rx_data_114),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_115(w_hssi_rx_pld_pcs_interface_pld_rx_data_115),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_116(w_hssi_rx_pld_pcs_interface_pld_rx_data_116),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_117(w_hssi_rx_pld_pcs_interface_pld_rx_data_117),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_118(w_hssi_rx_pld_pcs_interface_pld_rx_data_118),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_119(w_hssi_rx_pld_pcs_interface_pld_rx_data_119),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_120(w_hssi_rx_pld_pcs_interface_pld_rx_data_120),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_121(w_hssi_rx_pld_pcs_interface_pld_rx_data_121),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_122(w_hssi_rx_pld_pcs_interface_pld_rx_data_122),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_123(w_hssi_rx_pld_pcs_interface_pld_rx_data_123),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_124(w_hssi_rx_pld_pcs_interface_pld_rx_data_124),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_125(w_hssi_rx_pld_pcs_interface_pld_rx_data_125),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_126(w_hssi_rx_pld_pcs_interface_pld_rx_data_126),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_127(w_hssi_rx_pld_pcs_interface_pld_rx_data_127),
	.pld_cal_done_0(pld_cal_done_0),
	.avmm_readdata_0(avmm_readdata_0),
	.avmm_readdata_1(avmm_readdata_1),
	.avmm_readdata_2(avmm_readdata_2),
	.avmm_readdata_3(avmm_readdata_3),
	.avmm_readdata_4(avmm_readdata_4),
	.avmm_readdata_5(avmm_readdata_5),
	.avmm_readdata_6(avmm_readdata_6),
	.avmm_readdata_7(avmm_readdata_7),
	.out_pld_pma_pfdmode_lock(w_hssi_common_pld_pcs_interface_pld_pma_pfdmode_lock),
	.out_pld_pma_rxpll_lock(w_hssi_common_pld_pcs_interface_pld_pma_rxpll_lock),
	.out_pld_pcs_tx_clk_out(tx_clkout[0]),
	.out_tx_p(tx_serial_data[0]),
	.avmm_waitrequest_0(avmm_waitrequest_0),
	.reset_out_stage_0(reset_out_stage_0),
	.reset_out_stage_1(reset_out_stage_1),
	.reconfig_read_0(reconfig_read_0),
	.rx_digitalreset_0(rx_digitalreset_0),
	.rx_std_wa_patternalign_0(rx_std_wa_patternalign_0),
	.rx_coreclkin_0(rx_coreclkin_0),
	.reconfig_clk_0(reconfig_clk_0),
	.reconfig_write_0(reconfig_write_0),
	.reconfig_address_0(reconfig_address_0),
	.reconfig_address_1(reconfig_address_1),
	.reconfig_address_2(reconfig_address_2),
	.reconfig_address_3(reconfig_address_3),
	.reconfig_address_4(reconfig_address_4),
	.reconfig_address_5(reconfig_address_5),
	.reconfig_address_6(reconfig_address_6),
	.reconfig_address_7(reconfig_address_7),
	.reconfig_address_8(reconfig_address_8),
	.reconfig_writedata_0(reconfig_writedata_0),
	.reconfig_writedata_1(reconfig_writedata_1),
	.reconfig_writedata_2(reconfig_writedata_2),
	.reconfig_writedata_3(reconfig_writedata_3),
	.reconfig_writedata_4(reconfig_writedata_4),
	.reconfig_writedata_5(reconfig_writedata_5),
	.reconfig_writedata_6(reconfig_writedata_6),
	.reconfig_writedata_7(reconfig_writedata_7),
	.rx_seriallpbken_0(rx_seriallpbken_0),
	.tx_digitalreset_0(tx_digitalreset_0),
	.tx_coreclkin_0(tx_coreclkin_0),
	.tx_parallel_data_0(tx_parallel_data_0),
	.tx_parallel_data_1(tx_parallel_data_1),
	.tx_parallel_data_2(tx_parallel_data_2),
	.tx_parallel_data_3(tx_parallel_data_3),
	.tx_parallel_data_4(tx_parallel_data_4),
	.tx_parallel_data_5(tx_parallel_data_5),
	.tx_parallel_data_6(tx_parallel_data_6),
	.tx_parallel_data_7(tx_parallel_data_7),
	.tx_datak(tx_datak),
	.unused_tx_parallel_data_0(unused_tx_parallel_data_0),
	.unused_tx_parallel_data_1(unused_tx_parallel_data_1),
	.unused_tx_parallel_data_2(unused_tx_parallel_data_2),
	.unused_tx_parallel_data_3(unused_tx_parallel_data_3),
	.unused_tx_parallel_data_4(unused_tx_parallel_data_4),
	.unused_tx_parallel_data_5(unused_tx_parallel_data_5),
	.unused_tx_parallel_data_6(unused_tx_parallel_data_6),
	.unused_tx_parallel_data_7(unused_tx_parallel_data_7),
	.unused_tx_parallel_data_8(unused_tx_parallel_data_8),
	.unused_tx_parallel_data_9(unused_tx_parallel_data_9),
	.unused_tx_parallel_data_10(unused_tx_parallel_data_10),
	.unused_tx_parallel_data_11(unused_tx_parallel_data_11),
	.unused_tx_parallel_data_12(unused_tx_parallel_data_12),
	.unused_tx_parallel_data_13(unused_tx_parallel_data_13),
	.unused_tx_parallel_data_14(unused_tx_parallel_data_14),
	.unused_tx_parallel_data_15(unused_tx_parallel_data_15),
	.unused_tx_parallel_data_16(unused_tx_parallel_data_16),
	.unused_tx_parallel_data_17(unused_tx_parallel_data_17),
	.unused_tx_parallel_data_18(unused_tx_parallel_data_18),
	.unused_tx_parallel_data_19(unused_tx_parallel_data_19),
	.unused_tx_parallel_data_20(unused_tx_parallel_data_20),
	.unused_tx_parallel_data_21(unused_tx_parallel_data_21),
	.unused_tx_parallel_data_22(unused_tx_parallel_data_22),
	.unused_tx_parallel_data_23(unused_tx_parallel_data_23),
	.unused_tx_parallel_data_24(unused_tx_parallel_data_24),
	.unused_tx_parallel_data_25(unused_tx_parallel_data_25),
	.unused_tx_parallel_data_26(unused_tx_parallel_data_26),
	.unused_tx_parallel_data_27(unused_tx_parallel_data_27),
	.unused_tx_parallel_data_28(unused_tx_parallel_data_28),
	.unused_tx_parallel_data_29(unused_tx_parallel_data_29),
	.unused_tx_parallel_data_30(unused_tx_parallel_data_30),
	.unused_tx_parallel_data_31(unused_tx_parallel_data_31),
	.unused_tx_parallel_data_32(unused_tx_parallel_data_32),
	.unused_tx_parallel_data_33(unused_tx_parallel_data_33),
	.unused_tx_parallel_data_34(unused_tx_parallel_data_34),
	.unused_tx_parallel_data_35(unused_tx_parallel_data_35),
	.unused_tx_parallel_data_36(unused_tx_parallel_data_36),
	.unused_tx_parallel_data_37(unused_tx_parallel_data_37),
	.unused_tx_parallel_data_38(unused_tx_parallel_data_38),
	.unused_tx_parallel_data_39(unused_tx_parallel_data_39),
	.unused_tx_parallel_data_40(unused_tx_parallel_data_40),
	.unused_tx_parallel_data_41(unused_tx_parallel_data_41),
	.unused_tx_parallel_data_42(unused_tx_parallel_data_42),
	.unused_tx_parallel_data_43(unused_tx_parallel_data_43),
	.unused_tx_parallel_data_44(unused_tx_parallel_data_44),
	.unused_tx_parallel_data_45(unused_tx_parallel_data_45),
	.unused_tx_parallel_data_46(unused_tx_parallel_data_46),
	.unused_tx_parallel_data_47(unused_tx_parallel_data_47),
	.unused_tx_parallel_data_48(unused_tx_parallel_data_48),
	.unused_tx_parallel_data_49(unused_tx_parallel_data_49),
	.unused_tx_parallel_data_50(unused_tx_parallel_data_50),
	.unused_tx_parallel_data_51(unused_tx_parallel_data_51),
	.unused_tx_parallel_data_52(unused_tx_parallel_data_52),
	.unused_tx_parallel_data_53(unused_tx_parallel_data_53),
	.unused_tx_parallel_data_54(unused_tx_parallel_data_54),
	.unused_tx_parallel_data_55(unused_tx_parallel_data_55),
	.unused_tx_parallel_data_56(unused_tx_parallel_data_56),
	.unused_tx_parallel_data_57(unused_tx_parallel_data_57),
	.unused_tx_parallel_data_58(unused_tx_parallel_data_58),
	.unused_tx_parallel_data_59(unused_tx_parallel_data_59),
	.unused_tx_parallel_data_60(unused_tx_parallel_data_60),
	.unused_tx_parallel_data_61(unused_tx_parallel_data_61),
	.unused_tx_parallel_data_62(unused_tx_parallel_data_62),
	.unused_tx_parallel_data_63(unused_tx_parallel_data_63),
	.unused_tx_parallel_data_64(unused_tx_parallel_data_64),
	.unused_tx_parallel_data_65(unused_tx_parallel_data_65),
	.unused_tx_parallel_data_66(unused_tx_parallel_data_66),
	.unused_tx_parallel_data_67(unused_tx_parallel_data_67),
	.unused_tx_parallel_data_68(unused_tx_parallel_data_68),
	.unused_tx_parallel_data_69(unused_tx_parallel_data_69),
	.unused_tx_parallel_data_70(unused_tx_parallel_data_70),
	.unused_tx_parallel_data_71(unused_tx_parallel_data_71),
	.unused_tx_parallel_data_72(unused_tx_parallel_data_72),
	.unused_tx_parallel_data_73(unused_tx_parallel_data_73),
	.unused_tx_parallel_data_74(unused_tx_parallel_data_74),
	.unused_tx_parallel_data_75(unused_tx_parallel_data_75),
	.unused_tx_parallel_data_76(unused_tx_parallel_data_76),
	.unused_tx_parallel_data_77(unused_tx_parallel_data_77),
	.unused_tx_parallel_data_78(unused_tx_parallel_data_78),
	.unused_tx_parallel_data_79(unused_tx_parallel_data_79),
	.unused_tx_parallel_data_80(unused_tx_parallel_data_80),
	.unused_tx_parallel_data_81(unused_tx_parallel_data_81),
	.unused_tx_parallel_data_82(unused_tx_parallel_data_82),
	.unused_tx_parallel_data_83(unused_tx_parallel_data_83),
	.unused_tx_parallel_data_84(unused_tx_parallel_data_84),
	.unused_tx_parallel_data_85(unused_tx_parallel_data_85),
	.unused_tx_parallel_data_86(unused_tx_parallel_data_86),
	.unused_tx_parallel_data_87(unused_tx_parallel_data_87),
	.unused_tx_parallel_data_88(unused_tx_parallel_data_88),
	.unused_tx_parallel_data_89(unused_tx_parallel_data_89),
	.unused_tx_parallel_data_90(unused_tx_parallel_data_90),
	.unused_tx_parallel_data_91(unused_tx_parallel_data_91),
	.unused_tx_parallel_data_92(unused_tx_parallel_data_92),
	.unused_tx_parallel_data_93(unused_tx_parallel_data_93),
	.unused_tx_parallel_data_94(unused_tx_parallel_data_94),
	.unused_tx_parallel_data_95(unused_tx_parallel_data_95),
	.unused_tx_parallel_data_96(unused_tx_parallel_data_96),
	.unused_tx_parallel_data_97(unused_tx_parallel_data_97),
	.unused_tx_parallel_data_98(unused_tx_parallel_data_98),
	.unused_tx_parallel_data_99(unused_tx_parallel_data_99),
	.unused_tx_parallel_data_100(unused_tx_parallel_data_100),
	.unused_tx_parallel_data_101(unused_tx_parallel_data_101),
	.unused_tx_parallel_data_102(unused_tx_parallel_data_102),
	.unused_tx_parallel_data_103(unused_tx_parallel_data_103),
	.unused_tx_parallel_data_104(unused_tx_parallel_data_104),
	.unused_tx_parallel_data_105(unused_tx_parallel_data_105),
	.unused_tx_parallel_data_106(unused_tx_parallel_data_106),
	.unused_tx_parallel_data_107(unused_tx_parallel_data_107),
	.unused_tx_parallel_data_108(unused_tx_parallel_data_108),
	.unused_tx_parallel_data_109(unused_tx_parallel_data_109),
	.unused_tx_parallel_data_110(unused_tx_parallel_data_110),
	.unused_tx_parallel_data_111(unused_tx_parallel_data_111),
	.unused_tx_parallel_data_112(unused_tx_parallel_data_112),
	.unused_tx_parallel_data_113(unused_tx_parallel_data_113),
	.unused_tx_parallel_data_114(unused_tx_parallel_data_114),
	.unused_tx_parallel_data_115(unused_tx_parallel_data_115),
	.unused_tx_parallel_data_116(unused_tx_parallel_data_116),
	.unused_tx_parallel_data_117(unused_tx_parallel_data_117),
	.unused_tx_parallel_data_118(unused_tx_parallel_data_118),
	.rx_serial_data_0(rx_serial_data_0),
	.tx_serial_clk0_0(tx_serial_clk0_0),
	.rx_cdr_refclk0(rx_cdr_refclk0),
	.reconfig_reset_0(reconfig_reset_0));

endmodule

module wr_arria10_e3p1_det_phy_twentynm_xcvr_native (
	out_pld_pcs_rx_clk_out,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_0,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_1,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_2,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_3,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_5,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_6,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_7,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_8,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_9,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_10,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_11,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_12,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_13,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_14,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_15,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_16,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_17,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_18,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_19,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_20,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_21,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_22,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_23,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_24,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_25,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_26,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_27,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_28,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_29,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_30,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_31,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_32,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_33,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_34,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_35,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_36,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_37,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_38,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_39,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_40,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_41,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_42,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_43,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_44,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_45,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_46,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_47,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_48,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_49,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_50,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_51,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_52,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_53,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_54,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_55,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_56,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_57,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_58,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_59,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_60,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_61,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_62,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_63,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_64,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_65,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_66,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_67,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_68,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_69,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_70,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_71,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_72,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_73,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_74,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_75,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_76,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_77,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_78,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_79,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_80,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_81,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_82,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_83,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_84,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_85,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_86,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_87,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_88,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_89,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_90,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_91,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_92,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_93,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_94,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_95,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_96,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_97,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_98,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_99,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_100,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_101,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_102,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_103,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_104,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_105,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_106,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_107,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_108,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_109,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_110,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_111,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_112,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_113,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_114,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_115,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_116,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_117,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_118,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_119,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_120,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_121,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_122,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_123,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_124,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_125,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_126,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_127,
	pld_cal_done_0,
	avmm_readdata_0,
	avmm_readdata_1,
	avmm_readdata_2,
	avmm_readdata_3,
	avmm_readdata_4,
	avmm_readdata_5,
	avmm_readdata_6,
	avmm_readdata_7,
	out_pld_pma_pfdmode_lock,
	out_pld_pma_rxpll_lock,
	out_pld_pcs_tx_clk_out,
	out_tx_p,
	avmm_waitrequest_0,
	reset_out_stage_0,
	reset_out_stage_1,
	reconfig_read_0,
	rx_digitalreset_0,
	rx_std_wa_patternalign_0,
	rx_coreclkin_0,
	reconfig_clk_0,
	reconfig_write_0,
	reconfig_address_0,
	reconfig_address_1,
	reconfig_address_2,
	reconfig_address_3,
	reconfig_address_4,
	reconfig_address_5,
	reconfig_address_6,
	reconfig_address_7,
	reconfig_address_8,
	reconfig_writedata_0,
	reconfig_writedata_1,
	reconfig_writedata_2,
	reconfig_writedata_3,
	reconfig_writedata_4,
	reconfig_writedata_5,
	reconfig_writedata_6,
	reconfig_writedata_7,
	rx_seriallpbken_0,
	tx_digitalreset_0,
	tx_coreclkin_0,
	tx_parallel_data_0,
	tx_parallel_data_1,
	tx_parallel_data_2,
	tx_parallel_data_3,
	tx_parallel_data_4,
	tx_parallel_data_5,
	tx_parallel_data_6,
	tx_parallel_data_7,
	tx_datak,
	unused_tx_parallel_data_0,
	unused_tx_parallel_data_1,
	unused_tx_parallel_data_2,
	unused_tx_parallel_data_3,
	unused_tx_parallel_data_4,
	unused_tx_parallel_data_5,
	unused_tx_parallel_data_6,
	unused_tx_parallel_data_7,
	unused_tx_parallel_data_8,
	unused_tx_parallel_data_9,
	unused_tx_parallel_data_10,
	unused_tx_parallel_data_11,
	unused_tx_parallel_data_12,
	unused_tx_parallel_data_13,
	unused_tx_parallel_data_14,
	unused_tx_parallel_data_15,
	unused_tx_parallel_data_16,
	unused_tx_parallel_data_17,
	unused_tx_parallel_data_18,
	unused_tx_parallel_data_19,
	unused_tx_parallel_data_20,
	unused_tx_parallel_data_21,
	unused_tx_parallel_data_22,
	unused_tx_parallel_data_23,
	unused_tx_parallel_data_24,
	unused_tx_parallel_data_25,
	unused_tx_parallel_data_26,
	unused_tx_parallel_data_27,
	unused_tx_parallel_data_28,
	unused_tx_parallel_data_29,
	unused_tx_parallel_data_30,
	unused_tx_parallel_data_31,
	unused_tx_parallel_data_32,
	unused_tx_parallel_data_33,
	unused_tx_parallel_data_34,
	unused_tx_parallel_data_35,
	unused_tx_parallel_data_36,
	unused_tx_parallel_data_37,
	unused_tx_parallel_data_38,
	unused_tx_parallel_data_39,
	unused_tx_parallel_data_40,
	unused_tx_parallel_data_41,
	unused_tx_parallel_data_42,
	unused_tx_parallel_data_43,
	unused_tx_parallel_data_44,
	unused_tx_parallel_data_45,
	unused_tx_parallel_data_46,
	unused_tx_parallel_data_47,
	unused_tx_parallel_data_48,
	unused_tx_parallel_data_49,
	unused_tx_parallel_data_50,
	unused_tx_parallel_data_51,
	unused_tx_parallel_data_52,
	unused_tx_parallel_data_53,
	unused_tx_parallel_data_54,
	unused_tx_parallel_data_55,
	unused_tx_parallel_data_56,
	unused_tx_parallel_data_57,
	unused_tx_parallel_data_58,
	unused_tx_parallel_data_59,
	unused_tx_parallel_data_60,
	unused_tx_parallel_data_61,
	unused_tx_parallel_data_62,
	unused_tx_parallel_data_63,
	unused_tx_parallel_data_64,
	unused_tx_parallel_data_65,
	unused_tx_parallel_data_66,
	unused_tx_parallel_data_67,
	unused_tx_parallel_data_68,
	unused_tx_parallel_data_69,
	unused_tx_parallel_data_70,
	unused_tx_parallel_data_71,
	unused_tx_parallel_data_72,
	unused_tx_parallel_data_73,
	unused_tx_parallel_data_74,
	unused_tx_parallel_data_75,
	unused_tx_parallel_data_76,
	unused_tx_parallel_data_77,
	unused_tx_parallel_data_78,
	unused_tx_parallel_data_79,
	unused_tx_parallel_data_80,
	unused_tx_parallel_data_81,
	unused_tx_parallel_data_82,
	unused_tx_parallel_data_83,
	unused_tx_parallel_data_84,
	unused_tx_parallel_data_85,
	unused_tx_parallel_data_86,
	unused_tx_parallel_data_87,
	unused_tx_parallel_data_88,
	unused_tx_parallel_data_89,
	unused_tx_parallel_data_90,
	unused_tx_parallel_data_91,
	unused_tx_parallel_data_92,
	unused_tx_parallel_data_93,
	unused_tx_parallel_data_94,
	unused_tx_parallel_data_95,
	unused_tx_parallel_data_96,
	unused_tx_parallel_data_97,
	unused_tx_parallel_data_98,
	unused_tx_parallel_data_99,
	unused_tx_parallel_data_100,
	unused_tx_parallel_data_101,
	unused_tx_parallel_data_102,
	unused_tx_parallel_data_103,
	unused_tx_parallel_data_104,
	unused_tx_parallel_data_105,
	unused_tx_parallel_data_106,
	unused_tx_parallel_data_107,
	unused_tx_parallel_data_108,
	unused_tx_parallel_data_109,
	unused_tx_parallel_data_110,
	unused_tx_parallel_data_111,
	unused_tx_parallel_data_112,
	unused_tx_parallel_data_113,
	unused_tx_parallel_data_114,
	unused_tx_parallel_data_115,
	unused_tx_parallel_data_116,
	unused_tx_parallel_data_117,
	unused_tx_parallel_data_118,
	rx_serial_data_0,
	tx_serial_clk0_0,
	rx_cdr_refclk0,
	reconfig_reset_0)/* synthesis synthesis_greybox=1 */;
output 	out_pld_pcs_rx_clk_out;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_0;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_1;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_2;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_3;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_5;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_6;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_7;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_8;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_9;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_10;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_11;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_12;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_13;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_14;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_15;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_16;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_17;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_18;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_19;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_20;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_21;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_22;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_23;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_24;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_25;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_26;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_27;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_28;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_29;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_30;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_31;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_32;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_33;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_34;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_35;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_36;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_37;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_38;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_39;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_40;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_41;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_42;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_43;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_44;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_45;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_46;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_47;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_48;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_49;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_50;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_51;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_52;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_53;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_54;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_55;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_56;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_57;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_58;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_59;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_60;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_61;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_62;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_63;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_64;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_65;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_66;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_67;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_68;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_69;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_70;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_71;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_72;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_73;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_74;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_75;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_76;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_77;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_78;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_79;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_80;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_81;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_82;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_83;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_84;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_85;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_86;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_87;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_88;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_89;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_90;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_91;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_92;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_93;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_94;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_95;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_96;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_97;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_98;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_99;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_100;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_101;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_102;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_103;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_104;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_105;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_106;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_107;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_108;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_109;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_110;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_111;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_112;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_113;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_114;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_115;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_116;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_117;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_118;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_119;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_120;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_121;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_122;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_123;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_124;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_125;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_126;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_127;
output 	pld_cal_done_0;
output 	avmm_readdata_0;
output 	avmm_readdata_1;
output 	avmm_readdata_2;
output 	avmm_readdata_3;
output 	avmm_readdata_4;
output 	avmm_readdata_5;
output 	avmm_readdata_6;
output 	avmm_readdata_7;
output 	out_pld_pma_pfdmode_lock;
output 	out_pld_pma_rxpll_lock;
output 	out_pld_pcs_tx_clk_out;
output 	out_tx_p;
output 	avmm_waitrequest_0;
input 	reset_out_stage_0;
input 	reset_out_stage_1;
input 	reconfig_read_0;
input 	rx_digitalreset_0;
input 	rx_std_wa_patternalign_0;
input 	rx_coreclkin_0;
input 	reconfig_clk_0;
input 	reconfig_write_0;
input 	reconfig_address_0;
input 	reconfig_address_1;
input 	reconfig_address_2;
input 	reconfig_address_3;
input 	reconfig_address_4;
input 	reconfig_address_5;
input 	reconfig_address_6;
input 	reconfig_address_7;
input 	reconfig_address_8;
input 	reconfig_writedata_0;
input 	reconfig_writedata_1;
input 	reconfig_writedata_2;
input 	reconfig_writedata_3;
input 	reconfig_writedata_4;
input 	reconfig_writedata_5;
input 	reconfig_writedata_6;
input 	reconfig_writedata_7;
input 	rx_seriallpbken_0;
input 	tx_digitalreset_0;
input 	tx_coreclkin_0;
input 	tx_parallel_data_0;
input 	tx_parallel_data_1;
input 	tx_parallel_data_2;
input 	tx_parallel_data_3;
input 	tx_parallel_data_4;
input 	tx_parallel_data_5;
input 	tx_parallel_data_6;
input 	tx_parallel_data_7;
input 	tx_datak;
input 	unused_tx_parallel_data_0;
input 	unused_tx_parallel_data_1;
input 	unused_tx_parallel_data_2;
input 	unused_tx_parallel_data_3;
input 	unused_tx_parallel_data_4;
input 	unused_tx_parallel_data_5;
input 	unused_tx_parallel_data_6;
input 	unused_tx_parallel_data_7;
input 	unused_tx_parallel_data_8;
input 	unused_tx_parallel_data_9;
input 	unused_tx_parallel_data_10;
input 	unused_tx_parallel_data_11;
input 	unused_tx_parallel_data_12;
input 	unused_tx_parallel_data_13;
input 	unused_tx_parallel_data_14;
input 	unused_tx_parallel_data_15;
input 	unused_tx_parallel_data_16;
input 	unused_tx_parallel_data_17;
input 	unused_tx_parallel_data_18;
input 	unused_tx_parallel_data_19;
input 	unused_tx_parallel_data_20;
input 	unused_tx_parallel_data_21;
input 	unused_tx_parallel_data_22;
input 	unused_tx_parallel_data_23;
input 	unused_tx_parallel_data_24;
input 	unused_tx_parallel_data_25;
input 	unused_tx_parallel_data_26;
input 	unused_tx_parallel_data_27;
input 	unused_tx_parallel_data_28;
input 	unused_tx_parallel_data_29;
input 	unused_tx_parallel_data_30;
input 	unused_tx_parallel_data_31;
input 	unused_tx_parallel_data_32;
input 	unused_tx_parallel_data_33;
input 	unused_tx_parallel_data_34;
input 	unused_tx_parallel_data_35;
input 	unused_tx_parallel_data_36;
input 	unused_tx_parallel_data_37;
input 	unused_tx_parallel_data_38;
input 	unused_tx_parallel_data_39;
input 	unused_tx_parallel_data_40;
input 	unused_tx_parallel_data_41;
input 	unused_tx_parallel_data_42;
input 	unused_tx_parallel_data_43;
input 	unused_tx_parallel_data_44;
input 	unused_tx_parallel_data_45;
input 	unused_tx_parallel_data_46;
input 	unused_tx_parallel_data_47;
input 	unused_tx_parallel_data_48;
input 	unused_tx_parallel_data_49;
input 	unused_tx_parallel_data_50;
input 	unused_tx_parallel_data_51;
input 	unused_tx_parallel_data_52;
input 	unused_tx_parallel_data_53;
input 	unused_tx_parallel_data_54;
input 	unused_tx_parallel_data_55;
input 	unused_tx_parallel_data_56;
input 	unused_tx_parallel_data_57;
input 	unused_tx_parallel_data_58;
input 	unused_tx_parallel_data_59;
input 	unused_tx_parallel_data_60;
input 	unused_tx_parallel_data_61;
input 	unused_tx_parallel_data_62;
input 	unused_tx_parallel_data_63;
input 	unused_tx_parallel_data_64;
input 	unused_tx_parallel_data_65;
input 	unused_tx_parallel_data_66;
input 	unused_tx_parallel_data_67;
input 	unused_tx_parallel_data_68;
input 	unused_tx_parallel_data_69;
input 	unused_tx_parallel_data_70;
input 	unused_tx_parallel_data_71;
input 	unused_tx_parallel_data_72;
input 	unused_tx_parallel_data_73;
input 	unused_tx_parallel_data_74;
input 	unused_tx_parallel_data_75;
input 	unused_tx_parallel_data_76;
input 	unused_tx_parallel_data_77;
input 	unused_tx_parallel_data_78;
input 	unused_tx_parallel_data_79;
input 	unused_tx_parallel_data_80;
input 	unused_tx_parallel_data_81;
input 	unused_tx_parallel_data_82;
input 	unused_tx_parallel_data_83;
input 	unused_tx_parallel_data_84;
input 	unused_tx_parallel_data_85;
input 	unused_tx_parallel_data_86;
input 	unused_tx_parallel_data_87;
input 	unused_tx_parallel_data_88;
input 	unused_tx_parallel_data_89;
input 	unused_tx_parallel_data_90;
input 	unused_tx_parallel_data_91;
input 	unused_tx_parallel_data_92;
input 	unused_tx_parallel_data_93;
input 	unused_tx_parallel_data_94;
input 	unused_tx_parallel_data_95;
input 	unused_tx_parallel_data_96;
input 	unused_tx_parallel_data_97;
input 	unused_tx_parallel_data_98;
input 	unused_tx_parallel_data_99;
input 	unused_tx_parallel_data_100;
input 	unused_tx_parallel_data_101;
input 	unused_tx_parallel_data_102;
input 	unused_tx_parallel_data_103;
input 	unused_tx_parallel_data_104;
input 	unused_tx_parallel_data_105;
input 	unused_tx_parallel_data_106;
input 	unused_tx_parallel_data_107;
input 	unused_tx_parallel_data_108;
input 	unused_tx_parallel_data_109;
input 	unused_tx_parallel_data_110;
input 	unused_tx_parallel_data_111;
input 	unused_tx_parallel_data_112;
input 	unused_tx_parallel_data_113;
input 	unused_tx_parallel_data_114;
input 	unused_tx_parallel_data_115;
input 	unused_tx_parallel_data_116;
input 	unused_tx_parallel_data_117;
input 	unused_tx_parallel_data_118;
input 	rx_serial_data_0;
input 	tx_serial_clk0_0;
input 	rx_cdr_refclk0;
input 	reconfig_reset_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



wr_arria10_e3p1_det_phy_twentynm_xcvr_native_rev_20nm5 twentynm_xcvr_native_inst(
	.out_pld_pcs_rx_clk_out(out_pld_pcs_rx_clk_out),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3),
	.w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4(w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_0(w_hssi_rx_pld_pcs_interface_pld_rx_data_0),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_1(w_hssi_rx_pld_pcs_interface_pld_rx_data_1),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_2(w_hssi_rx_pld_pcs_interface_pld_rx_data_2),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_3(w_hssi_rx_pld_pcs_interface_pld_rx_data_3),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_4(w_hssi_rx_pld_pcs_interface_pld_rx_data_4),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_5(w_hssi_rx_pld_pcs_interface_pld_rx_data_5),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_6(w_hssi_rx_pld_pcs_interface_pld_rx_data_6),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_7(w_hssi_rx_pld_pcs_interface_pld_rx_data_7),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_8(w_hssi_rx_pld_pcs_interface_pld_rx_data_8),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_9(w_hssi_rx_pld_pcs_interface_pld_rx_data_9),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_10(w_hssi_rx_pld_pcs_interface_pld_rx_data_10),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_11(w_hssi_rx_pld_pcs_interface_pld_rx_data_11),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_12(w_hssi_rx_pld_pcs_interface_pld_rx_data_12),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_13(w_hssi_rx_pld_pcs_interface_pld_rx_data_13),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_14(w_hssi_rx_pld_pcs_interface_pld_rx_data_14),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_15(w_hssi_rx_pld_pcs_interface_pld_rx_data_15),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_16(w_hssi_rx_pld_pcs_interface_pld_rx_data_16),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_17(w_hssi_rx_pld_pcs_interface_pld_rx_data_17),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_18(w_hssi_rx_pld_pcs_interface_pld_rx_data_18),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_19(w_hssi_rx_pld_pcs_interface_pld_rx_data_19),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_20(w_hssi_rx_pld_pcs_interface_pld_rx_data_20),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_21(w_hssi_rx_pld_pcs_interface_pld_rx_data_21),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_22(w_hssi_rx_pld_pcs_interface_pld_rx_data_22),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_23(w_hssi_rx_pld_pcs_interface_pld_rx_data_23),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_24(w_hssi_rx_pld_pcs_interface_pld_rx_data_24),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_25(w_hssi_rx_pld_pcs_interface_pld_rx_data_25),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_26(w_hssi_rx_pld_pcs_interface_pld_rx_data_26),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_27(w_hssi_rx_pld_pcs_interface_pld_rx_data_27),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_28(w_hssi_rx_pld_pcs_interface_pld_rx_data_28),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_29(w_hssi_rx_pld_pcs_interface_pld_rx_data_29),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_30(w_hssi_rx_pld_pcs_interface_pld_rx_data_30),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_31(w_hssi_rx_pld_pcs_interface_pld_rx_data_31),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_32(w_hssi_rx_pld_pcs_interface_pld_rx_data_32),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_33(w_hssi_rx_pld_pcs_interface_pld_rx_data_33),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_34(w_hssi_rx_pld_pcs_interface_pld_rx_data_34),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_35(w_hssi_rx_pld_pcs_interface_pld_rx_data_35),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_36(w_hssi_rx_pld_pcs_interface_pld_rx_data_36),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_37(w_hssi_rx_pld_pcs_interface_pld_rx_data_37),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_38(w_hssi_rx_pld_pcs_interface_pld_rx_data_38),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_39(w_hssi_rx_pld_pcs_interface_pld_rx_data_39),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_40(w_hssi_rx_pld_pcs_interface_pld_rx_data_40),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_41(w_hssi_rx_pld_pcs_interface_pld_rx_data_41),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_42(w_hssi_rx_pld_pcs_interface_pld_rx_data_42),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_43(w_hssi_rx_pld_pcs_interface_pld_rx_data_43),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_44(w_hssi_rx_pld_pcs_interface_pld_rx_data_44),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_45(w_hssi_rx_pld_pcs_interface_pld_rx_data_45),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_46(w_hssi_rx_pld_pcs_interface_pld_rx_data_46),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_47(w_hssi_rx_pld_pcs_interface_pld_rx_data_47),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_48(w_hssi_rx_pld_pcs_interface_pld_rx_data_48),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_49(w_hssi_rx_pld_pcs_interface_pld_rx_data_49),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_50(w_hssi_rx_pld_pcs_interface_pld_rx_data_50),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_51(w_hssi_rx_pld_pcs_interface_pld_rx_data_51),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_52(w_hssi_rx_pld_pcs_interface_pld_rx_data_52),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_53(w_hssi_rx_pld_pcs_interface_pld_rx_data_53),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_54(w_hssi_rx_pld_pcs_interface_pld_rx_data_54),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_55(w_hssi_rx_pld_pcs_interface_pld_rx_data_55),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_56(w_hssi_rx_pld_pcs_interface_pld_rx_data_56),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_57(w_hssi_rx_pld_pcs_interface_pld_rx_data_57),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_58(w_hssi_rx_pld_pcs_interface_pld_rx_data_58),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_59(w_hssi_rx_pld_pcs_interface_pld_rx_data_59),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_60(w_hssi_rx_pld_pcs_interface_pld_rx_data_60),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_61(w_hssi_rx_pld_pcs_interface_pld_rx_data_61),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_62(w_hssi_rx_pld_pcs_interface_pld_rx_data_62),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_63(w_hssi_rx_pld_pcs_interface_pld_rx_data_63),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_64(w_hssi_rx_pld_pcs_interface_pld_rx_data_64),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_65(w_hssi_rx_pld_pcs_interface_pld_rx_data_65),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_66(w_hssi_rx_pld_pcs_interface_pld_rx_data_66),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_67(w_hssi_rx_pld_pcs_interface_pld_rx_data_67),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_68(w_hssi_rx_pld_pcs_interface_pld_rx_data_68),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_69(w_hssi_rx_pld_pcs_interface_pld_rx_data_69),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_70(w_hssi_rx_pld_pcs_interface_pld_rx_data_70),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_71(w_hssi_rx_pld_pcs_interface_pld_rx_data_71),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_72(w_hssi_rx_pld_pcs_interface_pld_rx_data_72),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_73(w_hssi_rx_pld_pcs_interface_pld_rx_data_73),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_74(w_hssi_rx_pld_pcs_interface_pld_rx_data_74),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_75(w_hssi_rx_pld_pcs_interface_pld_rx_data_75),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_76(w_hssi_rx_pld_pcs_interface_pld_rx_data_76),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_77(w_hssi_rx_pld_pcs_interface_pld_rx_data_77),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_78(w_hssi_rx_pld_pcs_interface_pld_rx_data_78),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_79(w_hssi_rx_pld_pcs_interface_pld_rx_data_79),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_80(w_hssi_rx_pld_pcs_interface_pld_rx_data_80),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_81(w_hssi_rx_pld_pcs_interface_pld_rx_data_81),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_82(w_hssi_rx_pld_pcs_interface_pld_rx_data_82),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_83(w_hssi_rx_pld_pcs_interface_pld_rx_data_83),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_84(w_hssi_rx_pld_pcs_interface_pld_rx_data_84),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_85(w_hssi_rx_pld_pcs_interface_pld_rx_data_85),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_86(w_hssi_rx_pld_pcs_interface_pld_rx_data_86),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_87(w_hssi_rx_pld_pcs_interface_pld_rx_data_87),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_88(w_hssi_rx_pld_pcs_interface_pld_rx_data_88),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_89(w_hssi_rx_pld_pcs_interface_pld_rx_data_89),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_90(w_hssi_rx_pld_pcs_interface_pld_rx_data_90),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_91(w_hssi_rx_pld_pcs_interface_pld_rx_data_91),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_92(w_hssi_rx_pld_pcs_interface_pld_rx_data_92),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_93(w_hssi_rx_pld_pcs_interface_pld_rx_data_93),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_94(w_hssi_rx_pld_pcs_interface_pld_rx_data_94),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_95(w_hssi_rx_pld_pcs_interface_pld_rx_data_95),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_96(w_hssi_rx_pld_pcs_interface_pld_rx_data_96),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_97(w_hssi_rx_pld_pcs_interface_pld_rx_data_97),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_98(w_hssi_rx_pld_pcs_interface_pld_rx_data_98),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_99(w_hssi_rx_pld_pcs_interface_pld_rx_data_99),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_100(w_hssi_rx_pld_pcs_interface_pld_rx_data_100),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_101(w_hssi_rx_pld_pcs_interface_pld_rx_data_101),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_102(w_hssi_rx_pld_pcs_interface_pld_rx_data_102),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_103(w_hssi_rx_pld_pcs_interface_pld_rx_data_103),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_104(w_hssi_rx_pld_pcs_interface_pld_rx_data_104),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_105(w_hssi_rx_pld_pcs_interface_pld_rx_data_105),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_106(w_hssi_rx_pld_pcs_interface_pld_rx_data_106),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_107(w_hssi_rx_pld_pcs_interface_pld_rx_data_107),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_108(w_hssi_rx_pld_pcs_interface_pld_rx_data_108),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_109(w_hssi_rx_pld_pcs_interface_pld_rx_data_109),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_110(w_hssi_rx_pld_pcs_interface_pld_rx_data_110),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_111(w_hssi_rx_pld_pcs_interface_pld_rx_data_111),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_112(w_hssi_rx_pld_pcs_interface_pld_rx_data_112),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_113(w_hssi_rx_pld_pcs_interface_pld_rx_data_113),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_114(w_hssi_rx_pld_pcs_interface_pld_rx_data_114),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_115(w_hssi_rx_pld_pcs_interface_pld_rx_data_115),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_116(w_hssi_rx_pld_pcs_interface_pld_rx_data_116),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_117(w_hssi_rx_pld_pcs_interface_pld_rx_data_117),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_118(w_hssi_rx_pld_pcs_interface_pld_rx_data_118),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_119(w_hssi_rx_pld_pcs_interface_pld_rx_data_119),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_120(w_hssi_rx_pld_pcs_interface_pld_rx_data_120),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_121(w_hssi_rx_pld_pcs_interface_pld_rx_data_121),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_122(w_hssi_rx_pld_pcs_interface_pld_rx_data_122),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_123(w_hssi_rx_pld_pcs_interface_pld_rx_data_123),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_124(w_hssi_rx_pld_pcs_interface_pld_rx_data_124),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_125(w_hssi_rx_pld_pcs_interface_pld_rx_data_125),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_126(w_hssi_rx_pld_pcs_interface_pld_rx_data_126),
	.w_hssi_rx_pld_pcs_interface_pld_rx_data_127(w_hssi_rx_pld_pcs_interface_pld_rx_data_127),
	.pld_cal_done_0(pld_cal_done_0),
	.avmm_readdata_0(avmm_readdata_0),
	.avmm_readdata_1(avmm_readdata_1),
	.avmm_readdata_2(avmm_readdata_2),
	.avmm_readdata_3(avmm_readdata_3),
	.avmm_readdata_4(avmm_readdata_4),
	.avmm_readdata_5(avmm_readdata_5),
	.avmm_readdata_6(avmm_readdata_6),
	.avmm_readdata_7(avmm_readdata_7),
	.out_pld_pma_pfdmode_lock(out_pld_pma_pfdmode_lock),
	.out_pld_pma_rxpll_lock(out_pld_pma_rxpll_lock),
	.out_pld_pcs_tx_clk_out(out_pld_pcs_tx_clk_out),
	.out_tx_p(out_tx_p),
	.avmm_waitrequest_0(avmm_waitrequest_0),
	.reset_out_stage_0(reset_out_stage_0),
	.reset_out_stage_1(reset_out_stage_1),
	.reconfig_read_0(reconfig_read_0),
	.rx_digitalreset_0(rx_digitalreset_0),
	.rx_std_wa_patternalign_0(rx_std_wa_patternalign_0),
	.rx_coreclkin_0(rx_coreclkin_0),
	.reconfig_clk_0(reconfig_clk_0),
	.reconfig_write_0(reconfig_write_0),
	.reconfig_address_0(reconfig_address_0),
	.reconfig_address_1(reconfig_address_1),
	.reconfig_address_2(reconfig_address_2),
	.reconfig_address_3(reconfig_address_3),
	.reconfig_address_4(reconfig_address_4),
	.reconfig_address_5(reconfig_address_5),
	.reconfig_address_6(reconfig_address_6),
	.reconfig_address_7(reconfig_address_7),
	.reconfig_address_8(reconfig_address_8),
	.reconfig_writedata_0(reconfig_writedata_0),
	.reconfig_writedata_1(reconfig_writedata_1),
	.reconfig_writedata_2(reconfig_writedata_2),
	.reconfig_writedata_3(reconfig_writedata_3),
	.reconfig_writedata_4(reconfig_writedata_4),
	.reconfig_writedata_5(reconfig_writedata_5),
	.reconfig_writedata_6(reconfig_writedata_6),
	.reconfig_writedata_7(reconfig_writedata_7),
	.rx_seriallpbken_0(rx_seriallpbken_0),
	.tx_digitalreset_0(tx_digitalreset_0),
	.tx_coreclkin_0(tx_coreclkin_0),
	.tx_parallel_data_0(tx_parallel_data_0),
	.tx_parallel_data_1(tx_parallel_data_1),
	.tx_parallel_data_2(tx_parallel_data_2),
	.tx_parallel_data_3(tx_parallel_data_3),
	.tx_parallel_data_4(tx_parallel_data_4),
	.tx_parallel_data_5(tx_parallel_data_5),
	.tx_parallel_data_6(tx_parallel_data_6),
	.tx_parallel_data_7(tx_parallel_data_7),
	.tx_datak(tx_datak),
	.unused_tx_parallel_data_0(unused_tx_parallel_data_0),
	.unused_tx_parallel_data_1(unused_tx_parallel_data_1),
	.unused_tx_parallel_data_2(unused_tx_parallel_data_2),
	.unused_tx_parallel_data_3(unused_tx_parallel_data_3),
	.unused_tx_parallel_data_4(unused_tx_parallel_data_4),
	.unused_tx_parallel_data_5(unused_tx_parallel_data_5),
	.unused_tx_parallel_data_6(unused_tx_parallel_data_6),
	.unused_tx_parallel_data_7(unused_tx_parallel_data_7),
	.unused_tx_parallel_data_8(unused_tx_parallel_data_8),
	.unused_tx_parallel_data_9(unused_tx_parallel_data_9),
	.unused_tx_parallel_data_10(unused_tx_parallel_data_10),
	.unused_tx_parallel_data_11(unused_tx_parallel_data_11),
	.unused_tx_parallel_data_12(unused_tx_parallel_data_12),
	.unused_tx_parallel_data_13(unused_tx_parallel_data_13),
	.unused_tx_parallel_data_14(unused_tx_parallel_data_14),
	.unused_tx_parallel_data_15(unused_tx_parallel_data_15),
	.unused_tx_parallel_data_16(unused_tx_parallel_data_16),
	.unused_tx_parallel_data_17(unused_tx_parallel_data_17),
	.unused_tx_parallel_data_18(unused_tx_parallel_data_18),
	.unused_tx_parallel_data_19(unused_tx_parallel_data_19),
	.unused_tx_parallel_data_20(unused_tx_parallel_data_20),
	.unused_tx_parallel_data_21(unused_tx_parallel_data_21),
	.unused_tx_parallel_data_22(unused_tx_parallel_data_22),
	.unused_tx_parallel_data_23(unused_tx_parallel_data_23),
	.unused_tx_parallel_data_24(unused_tx_parallel_data_24),
	.unused_tx_parallel_data_25(unused_tx_parallel_data_25),
	.unused_tx_parallel_data_26(unused_tx_parallel_data_26),
	.unused_tx_parallel_data_27(unused_tx_parallel_data_27),
	.unused_tx_parallel_data_28(unused_tx_parallel_data_28),
	.unused_tx_parallel_data_29(unused_tx_parallel_data_29),
	.unused_tx_parallel_data_30(unused_tx_parallel_data_30),
	.unused_tx_parallel_data_31(unused_tx_parallel_data_31),
	.unused_tx_parallel_data_32(unused_tx_parallel_data_32),
	.unused_tx_parallel_data_33(unused_tx_parallel_data_33),
	.unused_tx_parallel_data_34(unused_tx_parallel_data_34),
	.unused_tx_parallel_data_35(unused_tx_parallel_data_35),
	.unused_tx_parallel_data_36(unused_tx_parallel_data_36),
	.unused_tx_parallel_data_37(unused_tx_parallel_data_37),
	.unused_tx_parallel_data_38(unused_tx_parallel_data_38),
	.unused_tx_parallel_data_39(unused_tx_parallel_data_39),
	.unused_tx_parallel_data_40(unused_tx_parallel_data_40),
	.unused_tx_parallel_data_41(unused_tx_parallel_data_41),
	.unused_tx_parallel_data_42(unused_tx_parallel_data_42),
	.unused_tx_parallel_data_43(unused_tx_parallel_data_43),
	.unused_tx_parallel_data_44(unused_tx_parallel_data_44),
	.unused_tx_parallel_data_45(unused_tx_parallel_data_45),
	.unused_tx_parallel_data_46(unused_tx_parallel_data_46),
	.unused_tx_parallel_data_47(unused_tx_parallel_data_47),
	.unused_tx_parallel_data_48(unused_tx_parallel_data_48),
	.unused_tx_parallel_data_49(unused_tx_parallel_data_49),
	.unused_tx_parallel_data_50(unused_tx_parallel_data_50),
	.unused_tx_parallel_data_51(unused_tx_parallel_data_51),
	.unused_tx_parallel_data_52(unused_tx_parallel_data_52),
	.unused_tx_parallel_data_53(unused_tx_parallel_data_53),
	.unused_tx_parallel_data_54(unused_tx_parallel_data_54),
	.unused_tx_parallel_data_55(unused_tx_parallel_data_55),
	.unused_tx_parallel_data_56(unused_tx_parallel_data_56),
	.unused_tx_parallel_data_57(unused_tx_parallel_data_57),
	.unused_tx_parallel_data_58(unused_tx_parallel_data_58),
	.unused_tx_parallel_data_59(unused_tx_parallel_data_59),
	.unused_tx_parallel_data_60(unused_tx_parallel_data_60),
	.unused_tx_parallel_data_61(unused_tx_parallel_data_61),
	.unused_tx_parallel_data_62(unused_tx_parallel_data_62),
	.unused_tx_parallel_data_63(unused_tx_parallel_data_63),
	.unused_tx_parallel_data_64(unused_tx_parallel_data_64),
	.unused_tx_parallel_data_65(unused_tx_parallel_data_65),
	.unused_tx_parallel_data_66(unused_tx_parallel_data_66),
	.unused_tx_parallel_data_67(unused_tx_parallel_data_67),
	.unused_tx_parallel_data_68(unused_tx_parallel_data_68),
	.unused_tx_parallel_data_69(unused_tx_parallel_data_69),
	.unused_tx_parallel_data_70(unused_tx_parallel_data_70),
	.unused_tx_parallel_data_71(unused_tx_parallel_data_71),
	.unused_tx_parallel_data_72(unused_tx_parallel_data_72),
	.unused_tx_parallel_data_73(unused_tx_parallel_data_73),
	.unused_tx_parallel_data_74(unused_tx_parallel_data_74),
	.unused_tx_parallel_data_75(unused_tx_parallel_data_75),
	.unused_tx_parallel_data_76(unused_tx_parallel_data_76),
	.unused_tx_parallel_data_77(unused_tx_parallel_data_77),
	.unused_tx_parallel_data_78(unused_tx_parallel_data_78),
	.unused_tx_parallel_data_79(unused_tx_parallel_data_79),
	.unused_tx_parallel_data_80(unused_tx_parallel_data_80),
	.unused_tx_parallel_data_81(unused_tx_parallel_data_81),
	.unused_tx_parallel_data_82(unused_tx_parallel_data_82),
	.unused_tx_parallel_data_83(unused_tx_parallel_data_83),
	.unused_tx_parallel_data_84(unused_tx_parallel_data_84),
	.unused_tx_parallel_data_85(unused_tx_parallel_data_85),
	.unused_tx_parallel_data_86(unused_tx_parallel_data_86),
	.unused_tx_parallel_data_87(unused_tx_parallel_data_87),
	.unused_tx_parallel_data_88(unused_tx_parallel_data_88),
	.unused_tx_parallel_data_89(unused_tx_parallel_data_89),
	.unused_tx_parallel_data_90(unused_tx_parallel_data_90),
	.unused_tx_parallel_data_91(unused_tx_parallel_data_91),
	.unused_tx_parallel_data_92(unused_tx_parallel_data_92),
	.unused_tx_parallel_data_93(unused_tx_parallel_data_93),
	.unused_tx_parallel_data_94(unused_tx_parallel_data_94),
	.unused_tx_parallel_data_95(unused_tx_parallel_data_95),
	.unused_tx_parallel_data_96(unused_tx_parallel_data_96),
	.unused_tx_parallel_data_97(unused_tx_parallel_data_97),
	.unused_tx_parallel_data_98(unused_tx_parallel_data_98),
	.unused_tx_parallel_data_99(unused_tx_parallel_data_99),
	.unused_tx_parallel_data_100(unused_tx_parallel_data_100),
	.unused_tx_parallel_data_101(unused_tx_parallel_data_101),
	.unused_tx_parallel_data_102(unused_tx_parallel_data_102),
	.unused_tx_parallel_data_103(unused_tx_parallel_data_103),
	.unused_tx_parallel_data_104(unused_tx_parallel_data_104),
	.unused_tx_parallel_data_105(unused_tx_parallel_data_105),
	.unused_tx_parallel_data_106(unused_tx_parallel_data_106),
	.unused_tx_parallel_data_107(unused_tx_parallel_data_107),
	.unused_tx_parallel_data_108(unused_tx_parallel_data_108),
	.unused_tx_parallel_data_109(unused_tx_parallel_data_109),
	.unused_tx_parallel_data_110(unused_tx_parallel_data_110),
	.unused_tx_parallel_data_111(unused_tx_parallel_data_111),
	.unused_tx_parallel_data_112(unused_tx_parallel_data_112),
	.unused_tx_parallel_data_113(unused_tx_parallel_data_113),
	.unused_tx_parallel_data_114(unused_tx_parallel_data_114),
	.unused_tx_parallel_data_115(unused_tx_parallel_data_115),
	.unused_tx_parallel_data_116(unused_tx_parallel_data_116),
	.unused_tx_parallel_data_117(unused_tx_parallel_data_117),
	.unused_tx_parallel_data_118(unused_tx_parallel_data_118),
	.rx_serial_data_0(rx_serial_data_0),
	.tx_serial_clk0_0(tx_serial_clk0_0),
	.rx_cdr_refclk0(rx_cdr_refclk0),
	.reconfig_reset_0(reconfig_reset_0));

endmodule

module wr_arria10_e3p1_det_phy_twentynm_xcvr_native_rev_20nm5 (
	out_pld_pcs_rx_clk_out,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3,
	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_0,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_1,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_2,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_3,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_4,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_5,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_6,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_7,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_8,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_9,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_10,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_11,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_12,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_13,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_14,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_15,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_16,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_17,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_18,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_19,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_20,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_21,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_22,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_23,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_24,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_25,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_26,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_27,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_28,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_29,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_30,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_31,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_32,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_33,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_34,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_35,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_36,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_37,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_38,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_39,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_40,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_41,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_42,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_43,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_44,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_45,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_46,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_47,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_48,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_49,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_50,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_51,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_52,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_53,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_54,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_55,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_56,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_57,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_58,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_59,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_60,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_61,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_62,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_63,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_64,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_65,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_66,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_67,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_68,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_69,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_70,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_71,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_72,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_73,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_74,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_75,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_76,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_77,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_78,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_79,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_80,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_81,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_82,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_83,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_84,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_85,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_86,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_87,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_88,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_89,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_90,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_91,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_92,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_93,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_94,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_95,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_96,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_97,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_98,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_99,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_100,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_101,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_102,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_103,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_104,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_105,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_106,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_107,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_108,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_109,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_110,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_111,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_112,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_113,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_114,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_115,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_116,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_117,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_118,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_119,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_120,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_121,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_122,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_123,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_124,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_125,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_126,
	w_hssi_rx_pld_pcs_interface_pld_rx_data_127,
	pld_cal_done_0,
	avmm_readdata_0,
	avmm_readdata_1,
	avmm_readdata_2,
	avmm_readdata_3,
	avmm_readdata_4,
	avmm_readdata_5,
	avmm_readdata_6,
	avmm_readdata_7,
	out_pld_pma_pfdmode_lock,
	out_pld_pma_rxpll_lock,
	out_pld_pcs_tx_clk_out,
	out_tx_p,
	avmm_waitrequest_0,
	reset_out_stage_0,
	reset_out_stage_1,
	reconfig_read_0,
	rx_digitalreset_0,
	rx_std_wa_patternalign_0,
	rx_coreclkin_0,
	reconfig_clk_0,
	reconfig_write_0,
	reconfig_address_0,
	reconfig_address_1,
	reconfig_address_2,
	reconfig_address_3,
	reconfig_address_4,
	reconfig_address_5,
	reconfig_address_6,
	reconfig_address_7,
	reconfig_address_8,
	reconfig_writedata_0,
	reconfig_writedata_1,
	reconfig_writedata_2,
	reconfig_writedata_3,
	reconfig_writedata_4,
	reconfig_writedata_5,
	reconfig_writedata_6,
	reconfig_writedata_7,
	rx_seriallpbken_0,
	tx_digitalreset_0,
	tx_coreclkin_0,
	tx_parallel_data_0,
	tx_parallel_data_1,
	tx_parallel_data_2,
	tx_parallel_data_3,
	tx_parallel_data_4,
	tx_parallel_data_5,
	tx_parallel_data_6,
	tx_parallel_data_7,
	tx_datak,
	unused_tx_parallel_data_0,
	unused_tx_parallel_data_1,
	unused_tx_parallel_data_2,
	unused_tx_parallel_data_3,
	unused_tx_parallel_data_4,
	unused_tx_parallel_data_5,
	unused_tx_parallel_data_6,
	unused_tx_parallel_data_7,
	unused_tx_parallel_data_8,
	unused_tx_parallel_data_9,
	unused_tx_parallel_data_10,
	unused_tx_parallel_data_11,
	unused_tx_parallel_data_12,
	unused_tx_parallel_data_13,
	unused_tx_parallel_data_14,
	unused_tx_parallel_data_15,
	unused_tx_parallel_data_16,
	unused_tx_parallel_data_17,
	unused_tx_parallel_data_18,
	unused_tx_parallel_data_19,
	unused_tx_parallel_data_20,
	unused_tx_parallel_data_21,
	unused_tx_parallel_data_22,
	unused_tx_parallel_data_23,
	unused_tx_parallel_data_24,
	unused_tx_parallel_data_25,
	unused_tx_parallel_data_26,
	unused_tx_parallel_data_27,
	unused_tx_parallel_data_28,
	unused_tx_parallel_data_29,
	unused_tx_parallel_data_30,
	unused_tx_parallel_data_31,
	unused_tx_parallel_data_32,
	unused_tx_parallel_data_33,
	unused_tx_parallel_data_34,
	unused_tx_parallel_data_35,
	unused_tx_parallel_data_36,
	unused_tx_parallel_data_37,
	unused_tx_parallel_data_38,
	unused_tx_parallel_data_39,
	unused_tx_parallel_data_40,
	unused_tx_parallel_data_41,
	unused_tx_parallel_data_42,
	unused_tx_parallel_data_43,
	unused_tx_parallel_data_44,
	unused_tx_parallel_data_45,
	unused_tx_parallel_data_46,
	unused_tx_parallel_data_47,
	unused_tx_parallel_data_48,
	unused_tx_parallel_data_49,
	unused_tx_parallel_data_50,
	unused_tx_parallel_data_51,
	unused_tx_parallel_data_52,
	unused_tx_parallel_data_53,
	unused_tx_parallel_data_54,
	unused_tx_parallel_data_55,
	unused_tx_parallel_data_56,
	unused_tx_parallel_data_57,
	unused_tx_parallel_data_58,
	unused_tx_parallel_data_59,
	unused_tx_parallel_data_60,
	unused_tx_parallel_data_61,
	unused_tx_parallel_data_62,
	unused_tx_parallel_data_63,
	unused_tx_parallel_data_64,
	unused_tx_parallel_data_65,
	unused_tx_parallel_data_66,
	unused_tx_parallel_data_67,
	unused_tx_parallel_data_68,
	unused_tx_parallel_data_69,
	unused_tx_parallel_data_70,
	unused_tx_parallel_data_71,
	unused_tx_parallel_data_72,
	unused_tx_parallel_data_73,
	unused_tx_parallel_data_74,
	unused_tx_parallel_data_75,
	unused_tx_parallel_data_76,
	unused_tx_parallel_data_77,
	unused_tx_parallel_data_78,
	unused_tx_parallel_data_79,
	unused_tx_parallel_data_80,
	unused_tx_parallel_data_81,
	unused_tx_parallel_data_82,
	unused_tx_parallel_data_83,
	unused_tx_parallel_data_84,
	unused_tx_parallel_data_85,
	unused_tx_parallel_data_86,
	unused_tx_parallel_data_87,
	unused_tx_parallel_data_88,
	unused_tx_parallel_data_89,
	unused_tx_parallel_data_90,
	unused_tx_parallel_data_91,
	unused_tx_parallel_data_92,
	unused_tx_parallel_data_93,
	unused_tx_parallel_data_94,
	unused_tx_parallel_data_95,
	unused_tx_parallel_data_96,
	unused_tx_parallel_data_97,
	unused_tx_parallel_data_98,
	unused_tx_parallel_data_99,
	unused_tx_parallel_data_100,
	unused_tx_parallel_data_101,
	unused_tx_parallel_data_102,
	unused_tx_parallel_data_103,
	unused_tx_parallel_data_104,
	unused_tx_parallel_data_105,
	unused_tx_parallel_data_106,
	unused_tx_parallel_data_107,
	unused_tx_parallel_data_108,
	unused_tx_parallel_data_109,
	unused_tx_parallel_data_110,
	unused_tx_parallel_data_111,
	unused_tx_parallel_data_112,
	unused_tx_parallel_data_113,
	unused_tx_parallel_data_114,
	unused_tx_parallel_data_115,
	unused_tx_parallel_data_116,
	unused_tx_parallel_data_117,
	unused_tx_parallel_data_118,
	rx_serial_data_0,
	tx_serial_clk0_0,
	rx_cdr_refclk0,
	reconfig_reset_0)/* synthesis synthesis_greybox=1 */;
output 	out_pld_pcs_rx_clk_out;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3;
output 	w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_0;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_1;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_2;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_3;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_4;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_5;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_6;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_7;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_8;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_9;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_10;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_11;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_12;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_13;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_14;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_15;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_16;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_17;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_18;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_19;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_20;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_21;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_22;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_23;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_24;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_25;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_26;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_27;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_28;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_29;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_30;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_31;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_32;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_33;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_34;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_35;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_36;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_37;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_38;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_39;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_40;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_41;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_42;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_43;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_44;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_45;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_46;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_47;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_48;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_49;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_50;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_51;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_52;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_53;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_54;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_55;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_56;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_57;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_58;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_59;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_60;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_61;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_62;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_63;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_64;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_65;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_66;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_67;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_68;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_69;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_70;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_71;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_72;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_73;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_74;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_75;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_76;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_77;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_78;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_79;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_80;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_81;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_82;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_83;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_84;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_85;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_86;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_87;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_88;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_89;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_90;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_91;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_92;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_93;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_94;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_95;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_96;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_97;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_98;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_99;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_100;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_101;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_102;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_103;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_104;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_105;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_106;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_107;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_108;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_109;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_110;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_111;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_112;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_113;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_114;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_115;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_116;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_117;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_118;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_119;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_120;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_121;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_122;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_123;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_124;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_125;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_126;
output 	w_hssi_rx_pld_pcs_interface_pld_rx_data_127;
output 	pld_cal_done_0;
output 	avmm_readdata_0;
output 	avmm_readdata_1;
output 	avmm_readdata_2;
output 	avmm_readdata_3;
output 	avmm_readdata_4;
output 	avmm_readdata_5;
output 	avmm_readdata_6;
output 	avmm_readdata_7;
output 	out_pld_pma_pfdmode_lock;
output 	out_pld_pma_rxpll_lock;
output 	out_pld_pcs_tx_clk_out;
output 	out_tx_p;
output 	avmm_waitrequest_0;
input 	reset_out_stage_0;
input 	reset_out_stage_1;
input 	reconfig_read_0;
input 	rx_digitalreset_0;
input 	rx_std_wa_patternalign_0;
input 	rx_coreclkin_0;
input 	reconfig_clk_0;
input 	reconfig_write_0;
input 	reconfig_address_0;
input 	reconfig_address_1;
input 	reconfig_address_2;
input 	reconfig_address_3;
input 	reconfig_address_4;
input 	reconfig_address_5;
input 	reconfig_address_6;
input 	reconfig_address_7;
input 	reconfig_address_8;
input 	reconfig_writedata_0;
input 	reconfig_writedata_1;
input 	reconfig_writedata_2;
input 	reconfig_writedata_3;
input 	reconfig_writedata_4;
input 	reconfig_writedata_5;
input 	reconfig_writedata_6;
input 	reconfig_writedata_7;
input 	rx_seriallpbken_0;
input 	tx_digitalreset_0;
input 	tx_coreclkin_0;
input 	tx_parallel_data_0;
input 	tx_parallel_data_1;
input 	tx_parallel_data_2;
input 	tx_parallel_data_3;
input 	tx_parallel_data_4;
input 	tx_parallel_data_5;
input 	tx_parallel_data_6;
input 	tx_parallel_data_7;
input 	tx_datak;
input 	unused_tx_parallel_data_0;
input 	unused_tx_parallel_data_1;
input 	unused_tx_parallel_data_2;
input 	unused_tx_parallel_data_3;
input 	unused_tx_parallel_data_4;
input 	unused_tx_parallel_data_5;
input 	unused_tx_parallel_data_6;
input 	unused_tx_parallel_data_7;
input 	unused_tx_parallel_data_8;
input 	unused_tx_parallel_data_9;
input 	unused_tx_parallel_data_10;
input 	unused_tx_parallel_data_11;
input 	unused_tx_parallel_data_12;
input 	unused_tx_parallel_data_13;
input 	unused_tx_parallel_data_14;
input 	unused_tx_parallel_data_15;
input 	unused_tx_parallel_data_16;
input 	unused_tx_parallel_data_17;
input 	unused_tx_parallel_data_18;
input 	unused_tx_parallel_data_19;
input 	unused_tx_parallel_data_20;
input 	unused_tx_parallel_data_21;
input 	unused_tx_parallel_data_22;
input 	unused_tx_parallel_data_23;
input 	unused_tx_parallel_data_24;
input 	unused_tx_parallel_data_25;
input 	unused_tx_parallel_data_26;
input 	unused_tx_parallel_data_27;
input 	unused_tx_parallel_data_28;
input 	unused_tx_parallel_data_29;
input 	unused_tx_parallel_data_30;
input 	unused_tx_parallel_data_31;
input 	unused_tx_parallel_data_32;
input 	unused_tx_parallel_data_33;
input 	unused_tx_parallel_data_34;
input 	unused_tx_parallel_data_35;
input 	unused_tx_parallel_data_36;
input 	unused_tx_parallel_data_37;
input 	unused_tx_parallel_data_38;
input 	unused_tx_parallel_data_39;
input 	unused_tx_parallel_data_40;
input 	unused_tx_parallel_data_41;
input 	unused_tx_parallel_data_42;
input 	unused_tx_parallel_data_43;
input 	unused_tx_parallel_data_44;
input 	unused_tx_parallel_data_45;
input 	unused_tx_parallel_data_46;
input 	unused_tx_parallel_data_47;
input 	unused_tx_parallel_data_48;
input 	unused_tx_parallel_data_49;
input 	unused_tx_parallel_data_50;
input 	unused_tx_parallel_data_51;
input 	unused_tx_parallel_data_52;
input 	unused_tx_parallel_data_53;
input 	unused_tx_parallel_data_54;
input 	unused_tx_parallel_data_55;
input 	unused_tx_parallel_data_56;
input 	unused_tx_parallel_data_57;
input 	unused_tx_parallel_data_58;
input 	unused_tx_parallel_data_59;
input 	unused_tx_parallel_data_60;
input 	unused_tx_parallel_data_61;
input 	unused_tx_parallel_data_62;
input 	unused_tx_parallel_data_63;
input 	unused_tx_parallel_data_64;
input 	unused_tx_parallel_data_65;
input 	unused_tx_parallel_data_66;
input 	unused_tx_parallel_data_67;
input 	unused_tx_parallel_data_68;
input 	unused_tx_parallel_data_69;
input 	unused_tx_parallel_data_70;
input 	unused_tx_parallel_data_71;
input 	unused_tx_parallel_data_72;
input 	unused_tx_parallel_data_73;
input 	unused_tx_parallel_data_74;
input 	unused_tx_parallel_data_75;
input 	unused_tx_parallel_data_76;
input 	unused_tx_parallel_data_77;
input 	unused_tx_parallel_data_78;
input 	unused_tx_parallel_data_79;
input 	unused_tx_parallel_data_80;
input 	unused_tx_parallel_data_81;
input 	unused_tx_parallel_data_82;
input 	unused_tx_parallel_data_83;
input 	unused_tx_parallel_data_84;
input 	unused_tx_parallel_data_85;
input 	unused_tx_parallel_data_86;
input 	unused_tx_parallel_data_87;
input 	unused_tx_parallel_data_88;
input 	unused_tx_parallel_data_89;
input 	unused_tx_parallel_data_90;
input 	unused_tx_parallel_data_91;
input 	unused_tx_parallel_data_92;
input 	unused_tx_parallel_data_93;
input 	unused_tx_parallel_data_94;
input 	unused_tx_parallel_data_95;
input 	unused_tx_parallel_data_96;
input 	unused_tx_parallel_data_97;
input 	unused_tx_parallel_data_98;
input 	unused_tx_parallel_data_99;
input 	unused_tx_parallel_data_100;
input 	unused_tx_parallel_data_101;
input 	unused_tx_parallel_data_102;
input 	unused_tx_parallel_data_103;
input 	unused_tx_parallel_data_104;
input 	unused_tx_parallel_data_105;
input 	unused_tx_parallel_data_106;
input 	unused_tx_parallel_data_107;
input 	unused_tx_parallel_data_108;
input 	unused_tx_parallel_data_109;
input 	unused_tx_parallel_data_110;
input 	unused_tx_parallel_data_111;
input 	unused_tx_parallel_data_112;
input 	unused_tx_parallel_data_113;
input 	unused_tx_parallel_data_114;
input 	unused_tx_parallel_data_115;
input 	unused_tx_parallel_data_116;
input 	unused_tx_parallel_data_117;
input 	unused_tx_parallel_data_118;
input 	rx_serial_data_0;
input 	tx_serial_clk0_0;
input 	rx_cdr_refclk0;
input 	reconfig_reset_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[7] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_clk[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_read[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_rstn[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_write[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[1] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[2] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[3] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[4] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[5] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[6] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[7] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[8] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[0] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[1] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[2] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[3] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[4] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[5] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[6] ;
wire \inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[7] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_tx_buf_blockselect ;
wire \inst_twentynm_pma|w_pma_tx_buf_rx_detect_valid ;
wire \inst_twentynm_pma|w_pma_tx_buf_rx_found ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_blockselect ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rx_clkslip ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4] ;
wire \inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5] ;
wire \inst_twentynm_pma|w_pma_tx_ser_blockselect ;
wire \inst_twentynm_pma|w_pma_tx_ser_clk_divtx ;
wire \inst_twentynm_pma|w_pma_tx_ser_clk_divtx_user ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_cgb_blockselect ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_cgb_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_cgb_pcie_sw_done[0] ;
wire \inst_twentynm_pma|w_pma_cgb_pcie_sw_done[1] ;
wire \inst_twentynm_pma|w_pma_rx_deser_blockselect ;
wire \inst_twentynm_pma|w_pma_rx_deser_clkdiv ;
wire \inst_twentynm_pma|w_pma_rx_deser_clkdiv_user ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[0] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[1] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[2] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[3] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[4] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[5] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[6] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[7] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[8] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[9] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[10] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[11] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[12] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[13] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[14] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[15] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[16] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[17] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[18] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[19] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[20] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[21] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[22] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[23] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[24] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[25] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[26] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[27] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[28] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[29] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[30] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[31] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[32] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[33] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[34] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[35] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[36] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[37] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[38] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[39] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[40] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[41] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[42] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[43] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[44] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[45] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[46] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[47] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[48] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[49] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[50] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[51] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[52] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[53] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[54] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[55] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[56] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[57] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[58] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[59] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[60] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[61] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[62] ;
wire \inst_twentynm_pma|w_pma_rx_deser_dout[63] ;
wire \inst_twentynm_pma|w_pma_rx_buf_blockselect ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_rx_sd_blockselect ;
wire \inst_twentynm_pma|w_pma_rx_sd_sd ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_rx_odi_blockselect ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_blockselect ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_cdr_pll_blockselect ;
wire \inst_twentynm_pma|w_cdr_pll_clklow ;
wire \inst_twentynm_pma|w_cdr_pll_fref ;
wire \inst_twentynm_pma|w_cdr_pll_pfdmode_lock ;
wire \inst_twentynm_pma|w_cdr_pll_rxpll_lock ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_cdr_pll_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_blockselect ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[7] ;
wire \inst_twentynm_pma|w_pma_adapt_blockselect ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[0] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[1] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[2] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[3] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[4] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[5] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[6] ;
wire \inst_twentynm_pma|w_pma_adapt_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_blockselect ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_blockselect ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_early_eios ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltd_b ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltr ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ppm_lock ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bitslip ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[0] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[1] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[2] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[3] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[4] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[5] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[6] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[7] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[8] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[9] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[10] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[11] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[12] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[13] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[14] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[15] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[16] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[17] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[0] ;
wire \inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[1] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_blockselect ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_txpma_rstb ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[0] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[1] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[2] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[3] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[4] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[5] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[6] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[7] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62] ;
wire \inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63] ;


wr_arria10_e3p1_det_phy_twentynm_xcvr_avmm inst_twentynm_xcvr_avmm(
	.pcs_blockselect_rx_pcs_pld_if({\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_blockselect }),
	.pcs_avmmreaddata_rx_pcs_pld_if({\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[0] }),
	.chnl_pll_avmm_clk({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_clk[0] }),
	.pld_cal_done({pld_cal_done_0}),
	.chnl_pll_avmm_read({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_read[0] }),
	.chnl_pll_avmm_rstn({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_rstn[0] }),
	.chnl_pll_avmm_write({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_write[0] }),
	.avmm_readdata({avmm_readdata_7,avmm_readdata_6,avmm_readdata_5,avmm_readdata_4,avmm_readdata_3,avmm_readdata_2,avmm_readdata_1,avmm_readdata_0}),
	.chnl_pll_avmm_address({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[8] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[0] }),
	.chnl_pll_avmm_writedata({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[0] }),
	.pcs_blockselect_com_pcs_pld_if({\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_blockselect }),
	.pcs_avmmreaddata_com_pcs_pld_if({\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[5] ,
\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[4] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[2] ,
\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[0] }),
	.pcs_blockselect_tx_pcs_pld_if({\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_blockselect }),
	.pcs_avmmreaddata_tx_pcs_pld_if({\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[0] }),
	.pma_blockselect_tx_buf({\inst_twentynm_pma|w_pma_tx_buf_blockselect }),
	.pma_avmmreaddata_tx_buf({\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[0] }),
	.pcs_blockselect_10g_rx_pcs({\inst_twentynm_pcs|w_hssi_10g_rx_pcs_blockselect }),
	.pcs_avmmreaddata_10g_rx_pcs({\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_8g_rx_pcs({\inst_twentynm_pcs|w_hssi_8g_rx_pcs_blockselect }),
	.pcs_avmmreaddata_8g_rx_pcs({\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_pipe_gen1_2({\inst_twentynm_pcs|w_hssi_pipe_gen1_2_blockselect }),
	.pcs_avmmreaddata_pipe_gen1_2({\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[0] }),
	.pcs_blockselect_krfec_rx_pcs({\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_blockselect }),
	.pcs_avmmreaddata_krfec_rx_pcs({\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_rx_pcs_pma_if({\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_blockselect }),
	.pcs_avmmreaddata_rx_pcs_pma_if({\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[0] }),
	.pma_blockselect_tx_ser({\inst_twentynm_pma|w_pma_tx_ser_blockselect }),
	.pma_avmmreaddata_tx_ser({\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[0] }),
	.pma_blockselect_tx_cgb({\inst_twentynm_pma|w_pma_cgb_blockselect }),
	.pma_avmmreaddata_tx_cgb({\inst_twentynm_pma|w_pma_cgb_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_cgb_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[0] }),
	.pma_blockselect_rx_deser({\inst_twentynm_pma|w_pma_rx_deser_blockselect }),
	.pma_avmmreaddata_rx_deser({\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[0] }),
	.pma_blockselect_rx_buf({\inst_twentynm_pma|w_pma_rx_buf_blockselect }),
	.pma_avmmreaddata_rx_buf({\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[0] }),
	.pma_blockselect_rx_sd({\inst_twentynm_pma|w_pma_rx_sd_blockselect }),
	.pma_avmmreaddata_rx_sd({\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[0] }),
	.pma_blockselect_rx_odi({\inst_twentynm_pma|w_pma_rx_odi_blockselect }),
	.pma_avmmreaddata_rx_odi({\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[0] }),
	.pma_blockselect_rx_dfe({\inst_twentynm_pma|w_pma_rx_dfe_blockselect }),
	.pma_avmmreaddata_rx_dfe({\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[0] }),
	.pma_blockselect_cdr_pll({\inst_twentynm_pma|w_cdr_pll_blockselect }),
	.pma_avmmreaddata_cdr_pll({\inst_twentynm_pma|w_cdr_pll_avmmreaddata[7] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[6] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[5] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[4] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[3] ,
\inst_twentynm_pma|w_cdr_pll_avmmreaddata[2] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[1] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[0] }),
	.pma_blockselect_cdr_refclk_select({\inst_twentynm_pma|w_pma_cdr_refclk_blockselect }),
	.pma_avmmreaddata_cdr_refclk_select({\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[4] ,
\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[3] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[0] }),
	.pma_blockselect_pma_adapt({\inst_twentynm_pma|w_pma_adapt_blockselect }),
	.pma_avmmreaddata_pma_adapt({\inst_twentynm_pma|w_pma_adapt_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_adapt_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[0] }),
	.pcs_blockselect_8g_tx_pcs({\inst_twentynm_pcs|w_hssi_8g_tx_pcs_blockselect }),
	.pcs_avmmreaddata_8g_tx_pcs({\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_10g_tx_pcs({\inst_twentynm_pcs|w_hssi_10g_tx_pcs_blockselect }),
	.pcs_avmmreaddata_10g_tx_pcs({\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_gen3_rx_pcs({\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_blockselect }),
	.pcs_avmmreaddata_gen3_rx_pcs({\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_pipe_gen3({\inst_twentynm_pcs|w_hssi_pipe_gen3_blockselect }),
	.pcs_avmmreaddata_pipe_gen3({\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[0] }),
	.pcs_blockselect_gen3_tx_pcs({\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_blockselect }),
	.pcs_avmmreaddata_gen3_tx_pcs({\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_krfec_tx_pcs({\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_blockselect }),
	.pcs_avmmreaddata_krfec_tx_pcs({\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_fifo_rx_pcs({\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_blockselect }),
	.pcs_avmmreaddata_fifo_rx_pcs({\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_fifo_tx_pcs({\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_blockselect }),
	.pcs_avmmreaddata_fifo_tx_pcs({\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[0] }),
	.pcs_blockselect_com_pcs_pma_if({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_blockselect }),
	.pcs_avmmreaddata_com_pcs_pma_if({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[5] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[4] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[2] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[0] }),
	.pcs_blockselect_tx_pcs_pma_if({\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_blockselect }),
	.pcs_avmmreaddata_tx_pcs_pma_if({\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[0] }),
	.avmm_waitrequest_0(avmm_waitrequest_0),
	.avmm_read({reconfig_read_0}),
	.reconfig_clk_0(reconfig_clk_0),
	.avmm_write({reconfig_write_0}),
	.avmm_address({reconfig_address_8,reconfig_address_7,reconfig_address_6,reconfig_address_5,reconfig_address_4,reconfig_address_3,reconfig_address_2,reconfig_address_1,reconfig_address_0}),
	.avmm_writedata({reconfig_writedata_7,reconfig_writedata_6,reconfig_writedata_5,reconfig_writedata_4,reconfig_writedata_3,reconfig_writedata_2,reconfig_writedata_1,reconfig_writedata_0}),
	.reconfig_reset_0(reconfig_reset_0));

wr_arria10_e3p1_det_phy_twentynm_pcs_rev_20nm5 inst_twentynm_pcs(
	.out_blockselect_hssi_rx_pld_pcs_interface(\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_blockselect ),
	.out_pld_pcs_rx_clk_out(out_pld_pcs_rx_clk_out),
	.out_avmmreaddata_hssi_rx_pld_pcs_interface({\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_rx_pld_pcs_interface_avmmreaddata[0] }),
	.out_pld_8g_wa_boundary({w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_4,w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_3,w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_2,w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_1,w_hssi_rx_pld_pcs_interface_pld_8g_wa_boundary_0}),
	.out_pld_rx_data({w_hssi_rx_pld_pcs_interface_pld_rx_data_127,w_hssi_rx_pld_pcs_interface_pld_rx_data_126,w_hssi_rx_pld_pcs_interface_pld_rx_data_125,w_hssi_rx_pld_pcs_interface_pld_rx_data_124,w_hssi_rx_pld_pcs_interface_pld_rx_data_123,
w_hssi_rx_pld_pcs_interface_pld_rx_data_122,w_hssi_rx_pld_pcs_interface_pld_rx_data_121,w_hssi_rx_pld_pcs_interface_pld_rx_data_120,w_hssi_rx_pld_pcs_interface_pld_rx_data_119,w_hssi_rx_pld_pcs_interface_pld_rx_data_118,
w_hssi_rx_pld_pcs_interface_pld_rx_data_117,w_hssi_rx_pld_pcs_interface_pld_rx_data_116,w_hssi_rx_pld_pcs_interface_pld_rx_data_115,w_hssi_rx_pld_pcs_interface_pld_rx_data_114,w_hssi_rx_pld_pcs_interface_pld_rx_data_113,
w_hssi_rx_pld_pcs_interface_pld_rx_data_112,w_hssi_rx_pld_pcs_interface_pld_rx_data_111,w_hssi_rx_pld_pcs_interface_pld_rx_data_110,w_hssi_rx_pld_pcs_interface_pld_rx_data_109,w_hssi_rx_pld_pcs_interface_pld_rx_data_108,
w_hssi_rx_pld_pcs_interface_pld_rx_data_107,w_hssi_rx_pld_pcs_interface_pld_rx_data_106,w_hssi_rx_pld_pcs_interface_pld_rx_data_105,w_hssi_rx_pld_pcs_interface_pld_rx_data_104,w_hssi_rx_pld_pcs_interface_pld_rx_data_103,
w_hssi_rx_pld_pcs_interface_pld_rx_data_102,w_hssi_rx_pld_pcs_interface_pld_rx_data_101,w_hssi_rx_pld_pcs_interface_pld_rx_data_100,w_hssi_rx_pld_pcs_interface_pld_rx_data_99,w_hssi_rx_pld_pcs_interface_pld_rx_data_98,w_hssi_rx_pld_pcs_interface_pld_rx_data_97,
w_hssi_rx_pld_pcs_interface_pld_rx_data_96,w_hssi_rx_pld_pcs_interface_pld_rx_data_95,w_hssi_rx_pld_pcs_interface_pld_rx_data_94,w_hssi_rx_pld_pcs_interface_pld_rx_data_93,w_hssi_rx_pld_pcs_interface_pld_rx_data_92,w_hssi_rx_pld_pcs_interface_pld_rx_data_91,
w_hssi_rx_pld_pcs_interface_pld_rx_data_90,w_hssi_rx_pld_pcs_interface_pld_rx_data_89,w_hssi_rx_pld_pcs_interface_pld_rx_data_88,w_hssi_rx_pld_pcs_interface_pld_rx_data_87,w_hssi_rx_pld_pcs_interface_pld_rx_data_86,w_hssi_rx_pld_pcs_interface_pld_rx_data_85,
w_hssi_rx_pld_pcs_interface_pld_rx_data_84,w_hssi_rx_pld_pcs_interface_pld_rx_data_83,w_hssi_rx_pld_pcs_interface_pld_rx_data_82,w_hssi_rx_pld_pcs_interface_pld_rx_data_81,w_hssi_rx_pld_pcs_interface_pld_rx_data_80,w_hssi_rx_pld_pcs_interface_pld_rx_data_79,
w_hssi_rx_pld_pcs_interface_pld_rx_data_78,w_hssi_rx_pld_pcs_interface_pld_rx_data_77,w_hssi_rx_pld_pcs_interface_pld_rx_data_76,w_hssi_rx_pld_pcs_interface_pld_rx_data_75,w_hssi_rx_pld_pcs_interface_pld_rx_data_74,w_hssi_rx_pld_pcs_interface_pld_rx_data_73,
w_hssi_rx_pld_pcs_interface_pld_rx_data_72,w_hssi_rx_pld_pcs_interface_pld_rx_data_71,w_hssi_rx_pld_pcs_interface_pld_rx_data_70,w_hssi_rx_pld_pcs_interface_pld_rx_data_69,w_hssi_rx_pld_pcs_interface_pld_rx_data_68,w_hssi_rx_pld_pcs_interface_pld_rx_data_67,
w_hssi_rx_pld_pcs_interface_pld_rx_data_66,w_hssi_rx_pld_pcs_interface_pld_rx_data_65,w_hssi_rx_pld_pcs_interface_pld_rx_data_64,w_hssi_rx_pld_pcs_interface_pld_rx_data_63,w_hssi_rx_pld_pcs_interface_pld_rx_data_62,w_hssi_rx_pld_pcs_interface_pld_rx_data_61,
w_hssi_rx_pld_pcs_interface_pld_rx_data_60,w_hssi_rx_pld_pcs_interface_pld_rx_data_59,w_hssi_rx_pld_pcs_interface_pld_rx_data_58,w_hssi_rx_pld_pcs_interface_pld_rx_data_57,w_hssi_rx_pld_pcs_interface_pld_rx_data_56,w_hssi_rx_pld_pcs_interface_pld_rx_data_55,
w_hssi_rx_pld_pcs_interface_pld_rx_data_54,w_hssi_rx_pld_pcs_interface_pld_rx_data_53,w_hssi_rx_pld_pcs_interface_pld_rx_data_52,w_hssi_rx_pld_pcs_interface_pld_rx_data_51,w_hssi_rx_pld_pcs_interface_pld_rx_data_50,w_hssi_rx_pld_pcs_interface_pld_rx_data_49,
w_hssi_rx_pld_pcs_interface_pld_rx_data_48,w_hssi_rx_pld_pcs_interface_pld_rx_data_47,w_hssi_rx_pld_pcs_interface_pld_rx_data_46,w_hssi_rx_pld_pcs_interface_pld_rx_data_45,w_hssi_rx_pld_pcs_interface_pld_rx_data_44,w_hssi_rx_pld_pcs_interface_pld_rx_data_43,
w_hssi_rx_pld_pcs_interface_pld_rx_data_42,w_hssi_rx_pld_pcs_interface_pld_rx_data_41,w_hssi_rx_pld_pcs_interface_pld_rx_data_40,w_hssi_rx_pld_pcs_interface_pld_rx_data_39,w_hssi_rx_pld_pcs_interface_pld_rx_data_38,w_hssi_rx_pld_pcs_interface_pld_rx_data_37,
w_hssi_rx_pld_pcs_interface_pld_rx_data_36,w_hssi_rx_pld_pcs_interface_pld_rx_data_35,w_hssi_rx_pld_pcs_interface_pld_rx_data_34,w_hssi_rx_pld_pcs_interface_pld_rx_data_33,w_hssi_rx_pld_pcs_interface_pld_rx_data_32,w_hssi_rx_pld_pcs_interface_pld_rx_data_31,
w_hssi_rx_pld_pcs_interface_pld_rx_data_30,w_hssi_rx_pld_pcs_interface_pld_rx_data_29,w_hssi_rx_pld_pcs_interface_pld_rx_data_28,w_hssi_rx_pld_pcs_interface_pld_rx_data_27,w_hssi_rx_pld_pcs_interface_pld_rx_data_26,w_hssi_rx_pld_pcs_interface_pld_rx_data_25,
w_hssi_rx_pld_pcs_interface_pld_rx_data_24,w_hssi_rx_pld_pcs_interface_pld_rx_data_23,w_hssi_rx_pld_pcs_interface_pld_rx_data_22,w_hssi_rx_pld_pcs_interface_pld_rx_data_21,w_hssi_rx_pld_pcs_interface_pld_rx_data_20,w_hssi_rx_pld_pcs_interface_pld_rx_data_19,
w_hssi_rx_pld_pcs_interface_pld_rx_data_18,w_hssi_rx_pld_pcs_interface_pld_rx_data_17,w_hssi_rx_pld_pcs_interface_pld_rx_data_16,w_hssi_rx_pld_pcs_interface_pld_rx_data_15,w_hssi_rx_pld_pcs_interface_pld_rx_data_14,w_hssi_rx_pld_pcs_interface_pld_rx_data_13,
w_hssi_rx_pld_pcs_interface_pld_rx_data_12,w_hssi_rx_pld_pcs_interface_pld_rx_data_11,w_hssi_rx_pld_pcs_interface_pld_rx_data_10,w_hssi_rx_pld_pcs_interface_pld_rx_data_9,w_hssi_rx_pld_pcs_interface_pld_rx_data_8,w_hssi_rx_pld_pcs_interface_pld_rx_data_7,
w_hssi_rx_pld_pcs_interface_pld_rx_data_6,w_hssi_rx_pld_pcs_interface_pld_rx_data_5,w_hssi_rx_pld_pcs_interface_pld_rx_data_4,w_hssi_rx_pld_pcs_interface_pld_rx_data_3,w_hssi_rx_pld_pcs_interface_pld_rx_data_2,w_hssi_rx_pld_pcs_interface_pld_rx_data_1,
w_hssi_rx_pld_pcs_interface_pld_rx_data_0}),
	.in_avmmclk(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_clk[0] ),
	.in_avmmread(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_read[0] ),
	.in_avmmrstn(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_rstn[0] ),
	.in_avmmwrite(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_write[0] ),
	.in_avmmaddress({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[8] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[0] }),
	.in_avmmwritedata({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[0] }),
	.out_blockselect_hssi_common_pld_pcs_interface(\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_blockselect ),
	.out_pld_pma_pfdmode_lock(out_pld_pma_pfdmode_lock),
	.out_pld_pma_rxpll_lock(out_pld_pma_rxpll_lock),
	.out_avmmreaddata_hssi_common_pld_pcs_interface({\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[5] ,
\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[4] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[2] ,
\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_common_pld_pcs_interface_avmmreaddata[0] }),
	.out_blockselect_hssi_tx_pld_pcs_interface(\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_blockselect ),
	.out_pld_pcs_tx_clk_out(out_pld_pcs_tx_clk_out),
	.out_avmmreaddata_hssi_tx_pld_pcs_interface({\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_tx_pld_pcs_interface_avmmreaddata[0] }),
	.in_pma_rx_detect_valid(\inst_twentynm_pma|w_pma_tx_buf_rx_detect_valid ),
	.in_pma_rx_found(\inst_twentynm_pma|w_pma_tx_buf_rx_found ),
	.out_blockselect_hssi_10g_rx_pcs(\inst_twentynm_pcs|w_hssi_10g_rx_pcs_blockselect ),
	.out_avmmreaddata_hssi_10g_rx_pcs({\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_10g_rx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_8g_rx_pcs(\inst_twentynm_pcs|w_hssi_8g_rx_pcs_blockselect ),
	.out_avmmreaddata_hssi_8g_rx_pcs({\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_8g_rx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_pipe_gen1_2(\inst_twentynm_pcs|w_hssi_pipe_gen1_2_blockselect ),
	.out_avmmreaddata_hssi_pipe_gen1_2({\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_pipe_gen1_2_avmmreaddata[0] }),
	.out_blockselect_hssi_krfec_rx_pcs(\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_blockselect ),
	.out_avmmreaddata_hssi_krfec_rx_pcs({\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_krfec_rx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_rx_pcs_pma_interface(\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_blockselect ),
	.out_pma_rx_clkslip(\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rx_clkslip ),
	.out_pma_rxpma_rstb(\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb ),
	.out_avmmreaddata_hssi_rx_pcs_pma_interface({\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_avmmreaddata[0] }),
	.out_pma_eye_monitor({\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3] ,
\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0] }),
	.in_pma_tx_pma_clk(\inst_twentynm_pma|w_pma_tx_ser_clk_divtx ),
	.in_pma_tx_clkdiv_user(\inst_twentynm_pma|w_pma_tx_ser_clk_divtx_user ),
	.in_pma_pcie_sw_done({\inst_twentynm_pma|w_pma_cgb_pcie_sw_done[1] ,\inst_twentynm_pma|w_pma_cgb_pcie_sw_done[0] }),
	.in_pma_rx_pma_clk(\inst_twentynm_pma|w_pma_rx_deser_clkdiv ),
	.in_pma_rx_clkdiv_user(\inst_twentynm_pma|w_pma_rx_deser_clkdiv_user ),
	.in_pma_rx_pma_data({\inst_twentynm_pma|w_pma_rx_deser_dout[63] ,\inst_twentynm_pma|w_pma_rx_deser_dout[62] ,\inst_twentynm_pma|w_pma_rx_deser_dout[61] ,\inst_twentynm_pma|w_pma_rx_deser_dout[60] ,\inst_twentynm_pma|w_pma_rx_deser_dout[59] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[58] ,\inst_twentynm_pma|w_pma_rx_deser_dout[57] ,\inst_twentynm_pma|w_pma_rx_deser_dout[56] ,\inst_twentynm_pma|w_pma_rx_deser_dout[55] ,\inst_twentynm_pma|w_pma_rx_deser_dout[54] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[53] ,\inst_twentynm_pma|w_pma_rx_deser_dout[52] ,\inst_twentynm_pma|w_pma_rx_deser_dout[51] ,\inst_twentynm_pma|w_pma_rx_deser_dout[50] ,\inst_twentynm_pma|w_pma_rx_deser_dout[49] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[48] ,\inst_twentynm_pma|w_pma_rx_deser_dout[47] ,\inst_twentynm_pma|w_pma_rx_deser_dout[46] ,\inst_twentynm_pma|w_pma_rx_deser_dout[45] ,\inst_twentynm_pma|w_pma_rx_deser_dout[44] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[43] ,\inst_twentynm_pma|w_pma_rx_deser_dout[42] ,\inst_twentynm_pma|w_pma_rx_deser_dout[41] ,\inst_twentynm_pma|w_pma_rx_deser_dout[40] ,\inst_twentynm_pma|w_pma_rx_deser_dout[39] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[38] ,\inst_twentynm_pma|w_pma_rx_deser_dout[37] ,\inst_twentynm_pma|w_pma_rx_deser_dout[36] ,\inst_twentynm_pma|w_pma_rx_deser_dout[35] ,\inst_twentynm_pma|w_pma_rx_deser_dout[34] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[33] ,\inst_twentynm_pma|w_pma_rx_deser_dout[32] ,\inst_twentynm_pma|w_pma_rx_deser_dout[31] ,\inst_twentynm_pma|w_pma_rx_deser_dout[30] ,\inst_twentynm_pma|w_pma_rx_deser_dout[29] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[28] ,\inst_twentynm_pma|w_pma_rx_deser_dout[27] ,\inst_twentynm_pma|w_pma_rx_deser_dout[26] ,\inst_twentynm_pma|w_pma_rx_deser_dout[25] ,\inst_twentynm_pma|w_pma_rx_deser_dout[24] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[23] ,\inst_twentynm_pma|w_pma_rx_deser_dout[22] ,\inst_twentynm_pma|w_pma_rx_deser_dout[21] ,\inst_twentynm_pma|w_pma_rx_deser_dout[20] ,\inst_twentynm_pma|w_pma_rx_deser_dout[19] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[18] ,\inst_twentynm_pma|w_pma_rx_deser_dout[17] ,\inst_twentynm_pma|w_pma_rx_deser_dout[16] ,\inst_twentynm_pma|w_pma_rx_deser_dout[15] ,\inst_twentynm_pma|w_pma_rx_deser_dout[14] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[13] ,\inst_twentynm_pma|w_pma_rx_deser_dout[12] ,\inst_twentynm_pma|w_pma_rx_deser_dout[11] ,\inst_twentynm_pma|w_pma_rx_deser_dout[10] ,\inst_twentynm_pma|w_pma_rx_deser_dout[9] ,\inst_twentynm_pma|w_pma_rx_deser_dout[8] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[7] ,\inst_twentynm_pma|w_pma_rx_deser_dout[6] ,\inst_twentynm_pma|w_pma_rx_deser_dout[5] ,\inst_twentynm_pma|w_pma_rx_deser_dout[4] ,\inst_twentynm_pma|w_pma_rx_deser_dout[3] ,\inst_twentynm_pma|w_pma_rx_deser_dout[2] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[1] ,\inst_twentynm_pma|w_pma_rx_deser_dout[0] }),
	.in_pma_signal_det(\inst_twentynm_pma|w_pma_rx_sd_sd ),
	.in_pma_clklow(\inst_twentynm_pma|w_cdr_pll_clklow ),
	.in_pma_fref(\inst_twentynm_pma|w_cdr_pll_fref ),
	.in_pma_pfdmode_lock(\inst_twentynm_pma|w_cdr_pll_pfdmode_lock ),
	.in_pma_rxpll_lock(\inst_twentynm_pma|w_cdr_pll_rxpll_lock ),
	.out_blockselect_hssi_8g_tx_pcs(\inst_twentynm_pcs|w_hssi_8g_tx_pcs_blockselect ),
	.out_avmmreaddata_hssi_8g_tx_pcs({\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_8g_tx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_10g_tx_pcs(\inst_twentynm_pcs|w_hssi_10g_tx_pcs_blockselect ),
	.out_avmmreaddata_hssi_10g_tx_pcs({\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_10g_tx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_gen3_rx_pcs(\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_blockselect ),
	.out_avmmreaddata_hssi_gen3_rx_pcs({\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_gen3_rx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_pipe_gen3(\inst_twentynm_pcs|w_hssi_pipe_gen3_blockselect ),
	.out_avmmreaddata_hssi_pipe_gen3({\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_pipe_gen3_avmmreaddata[0] }),
	.out_blockselect_hssi_gen3_tx_pcs(\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_blockselect ),
	.out_avmmreaddata_hssi_gen3_tx_pcs({\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_gen3_tx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_krfec_tx_pcs(\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_blockselect ),
	.out_avmmreaddata_hssi_krfec_tx_pcs({\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_krfec_tx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_fifo_rx_pcs(\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_blockselect ),
	.out_avmmreaddata_hssi_fifo_rx_pcs({\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_fifo_rx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_fifo_tx_pcs(\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_blockselect ),
	.out_avmmreaddata_hssi_fifo_tx_pcs({\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_fifo_tx_pcs_avmmreaddata[0] }),
	.out_blockselect_hssi_common_pcs_pma_interface(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_blockselect ),
	.out_pma_early_eios(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_early_eios ),
	.out_pma_ltd_b(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltd_b ),
	.out_pma_ltr(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltr ),
	.out_pma_ppm_lock(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ppm_lock ),
	.out_pma_rs_lpbk_b(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b ),
	.out_pma_rx_qpi_pullup(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup ),
	.out_pma_tx_bitslip(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bitslip ),
	.out_pma_tx_bonding_rstb(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb ),
	.out_pma_tx_qpi_pulldn(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn ),
	.out_pma_tx_qpi_pullup(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup ),
	.out_pma_tx_txdetectrx(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx ),
	.out_avmmreaddata_hssi_common_pcs_pma_interface({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[5] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[4] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[2] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_avmmreaddata[0] }),
	.out_pma_current_coeff({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[17] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[16] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[15] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[14] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[13] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[12] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[11] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[10] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[9] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[8] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[7] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[6] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[5] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[4] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[3] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[2] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[0] }),
	.out_pma_pcie_switch({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[0] }),
	.out_blockselect_hssi_tx_pcs_pma_interface(\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_blockselect ),
	.out_pma_tx_elec_idle(\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle ),
	.out_pma_txpma_rstb(\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_txpma_rstb ),
	.out_avmmreaddata_hssi_tx_pcs_pma_interface({\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[7] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[6] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[5] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[4] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[3] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[2] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[1] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_avmmreaddata[0] }),
	.out_pma_tx_pma_data({\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0] }),
	.in_pld_pma_txpma_rstb(reset_out_stage_0),
	.in_pld_pma_rxpma_rstb(reset_out_stage_1),
	.in_pld_10g_krfec_rx_pld_rst_n(rx_digitalreset_0),
	.in_pld_8g_g3_rx_pld_rst_n(rx_digitalreset_0),
	.in_pld_pmaif_rx_pld_rst_n(rx_digitalreset_0),
	.in_pld_8g_encdt(rx_std_wa_patternalign_0),
	.in_pld_rx_clk(rx_coreclkin_0),
	.in_pld_pma_rs_lpbk_b(rx_seriallpbken_0),
	.in_pld_10g_krfec_tx_pld_rst_n(tx_digitalreset_0),
	.in_pld_8g_g3_tx_pld_rst_n(tx_digitalreset_0),
	.in_pld_pmaif_tx_pld_rst_n(tx_digitalreset_0),
	.in_pld_tx_clk(tx_coreclkin_0),
	.in_pld_tx_data({unused_tx_parallel_data_118,unused_tx_parallel_data_117,unused_tx_parallel_data_116,unused_tx_parallel_data_115,unused_tx_parallel_data_114,unused_tx_parallel_data_113,unused_tx_parallel_data_112,unused_tx_parallel_data_111,unused_tx_parallel_data_110,
unused_tx_parallel_data_109,unused_tx_parallel_data_108,unused_tx_parallel_data_107,unused_tx_parallel_data_106,unused_tx_parallel_data_105,unused_tx_parallel_data_104,unused_tx_parallel_data_103,unused_tx_parallel_data_102,unused_tx_parallel_data_101,
unused_tx_parallel_data_100,unused_tx_parallel_data_99,unused_tx_parallel_data_98,unused_tx_parallel_data_97,unused_tx_parallel_data_96,unused_tx_parallel_data_95,unused_tx_parallel_data_94,unused_tx_parallel_data_93,unused_tx_parallel_data_92,
unused_tx_parallel_data_91,unused_tx_parallel_data_90,unused_tx_parallel_data_89,unused_tx_parallel_data_88,unused_tx_parallel_data_87,unused_tx_parallel_data_86,unused_tx_parallel_data_85,unused_tx_parallel_data_84,unused_tx_parallel_data_83,
unused_tx_parallel_data_82,unused_tx_parallel_data_81,unused_tx_parallel_data_80,unused_tx_parallel_data_79,unused_tx_parallel_data_78,unused_tx_parallel_data_77,unused_tx_parallel_data_76,unused_tx_parallel_data_75,unused_tx_parallel_data_74,
unused_tx_parallel_data_73,unused_tx_parallel_data_72,unused_tx_parallel_data_71,unused_tx_parallel_data_70,unused_tx_parallel_data_69,unused_tx_parallel_data_68,unused_tx_parallel_data_67,unused_tx_parallel_data_66,unused_tx_parallel_data_65,
unused_tx_parallel_data_64,unused_tx_parallel_data_63,unused_tx_parallel_data_62,unused_tx_parallel_data_61,unused_tx_parallel_data_60,unused_tx_parallel_data_59,unused_tx_parallel_data_58,unused_tx_parallel_data_57,unused_tx_parallel_data_56,
unused_tx_parallel_data_55,unused_tx_parallel_data_54,unused_tx_parallel_data_53,unused_tx_parallel_data_52,unused_tx_parallel_data_51,unused_tx_parallel_data_50,unused_tx_parallel_data_49,unused_tx_parallel_data_48,unused_tx_parallel_data_47,
unused_tx_parallel_data_46,unused_tx_parallel_data_45,unused_tx_parallel_data_44,unused_tx_parallel_data_43,unused_tx_parallel_data_42,unused_tx_parallel_data_41,unused_tx_parallel_data_40,unused_tx_parallel_data_39,unused_tx_parallel_data_38,
unused_tx_parallel_data_37,unused_tx_parallel_data_36,unused_tx_parallel_data_35,unused_tx_parallel_data_34,unused_tx_parallel_data_33,unused_tx_parallel_data_32,unused_tx_parallel_data_31,unused_tx_parallel_data_30,unused_tx_parallel_data_29,
unused_tx_parallel_data_28,unused_tx_parallel_data_27,unused_tx_parallel_data_26,unused_tx_parallel_data_25,unused_tx_parallel_data_24,unused_tx_parallel_data_23,unused_tx_parallel_data_22,unused_tx_parallel_data_21,unused_tx_parallel_data_20,
unused_tx_parallel_data_19,unused_tx_parallel_data_18,unused_tx_parallel_data_17,unused_tx_parallel_data_16,unused_tx_parallel_data_15,unused_tx_parallel_data_14,unused_tx_parallel_data_13,unused_tx_parallel_data_12,unused_tx_parallel_data_11,
unused_tx_parallel_data_10,unused_tx_parallel_data_9,unused_tx_parallel_data_8,unused_tx_parallel_data_7,unused_tx_parallel_data_6,unused_tx_parallel_data_5,unused_tx_parallel_data_4,unused_tx_parallel_data_3,unused_tx_parallel_data_2,unused_tx_parallel_data_1,
unused_tx_parallel_data_0,tx_datak,tx_parallel_data_7,tx_parallel_data_6,tx_parallel_data_5,tx_parallel_data_4,tx_parallel_data_3,tx_parallel_data_2,tx_parallel_data_1,tx_parallel_data_0}));

wr_arria10_e3p1_det_phy_twentynm_pma_rev_20nm5 inst_twentynm_pma(
	.in_avmmclk(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_clk[0] ),
	.in_avmmread(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_read[0] ),
	.in_avmmrstn(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_rstn[0] ),
	.in_avmmwrite(\inst_twentynm_xcvr_avmm|chnl_pll_avmm_write[0] ),
	.in_avmmaddress({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[8] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_address[0] }),
	.in_avmmwritedata({\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[7] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[6] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[5] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[4] ,
\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[3] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[2] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[1] ,\inst_twentynm_xcvr_avmm|chnl_pll_avmm_writedata[0] }),
	.out_blockselect_pma_tx_buf(\inst_twentynm_pma|w_pma_tx_buf_blockselect ),
	.out_rx_detect_valid(\inst_twentynm_pma|w_pma_tx_buf_rx_detect_valid ),
	.out_rx_found(\inst_twentynm_pma|w_pma_tx_buf_rx_found ),
	.out_tx_p(out_tx_p),
	.out_avmmreaddata_pma_tx_buf({\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_tx_buf_avmmreaddata[0] }),
	.in_rx_bitslip(\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rx_clkslip ),
	.in_rx_pma_rstb(\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_rxpma_rstb ),
	.in_eye_monitor({\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[5] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[4] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[3] ,
\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[2] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[1] ,\inst_twentynm_pcs|w_hssi_rx_pcs_pma_interface_pma_eye_monitor[0] }),
	.out_blockselect_pma_tx_ser(\inst_twentynm_pma|w_pma_tx_ser_blockselect ),
	.out_iqtxrxclk_out1(\inst_twentynm_pma|w_pma_tx_ser_clk_divtx ),
	.out_clkdiv_tx_user(\inst_twentynm_pma|w_pma_tx_ser_clk_divtx_user ),
	.out_avmmreaddata_pma_tx_ser({\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_tx_ser_avmmreaddata[0] }),
	.out_blockselect_pma_cgb(\inst_twentynm_pma|w_pma_cgb_blockselect ),
	.out_avmmreaddata_pma_cgb({\inst_twentynm_pma|w_pma_cgb_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_cgb_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_cgb_avmmreaddata[0] }),
	.out_pcie_sw_done({\inst_twentynm_pma|w_pma_cgb_pcie_sw_done[1] ,\inst_twentynm_pma|w_pma_cgb_pcie_sw_done[0] }),
	.out_blockselect_pma_rx_deser(\inst_twentynm_pma|w_pma_rx_deser_blockselect ),
	.out_clkdiv_rx(\inst_twentynm_pma|w_pma_rx_deser_clkdiv ),
	.out_clkdiv_rx_user(\inst_twentynm_pma|w_pma_rx_deser_clkdiv_user ),
	.out_avmmreaddata_pma_rx_deser({\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_deser_avmmreaddata[0] }),
	.out_rxdata({\inst_twentynm_pma|w_pma_rx_deser_dout[63] ,\inst_twentynm_pma|w_pma_rx_deser_dout[62] ,\inst_twentynm_pma|w_pma_rx_deser_dout[61] ,\inst_twentynm_pma|w_pma_rx_deser_dout[60] ,\inst_twentynm_pma|w_pma_rx_deser_dout[59] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[58] ,\inst_twentynm_pma|w_pma_rx_deser_dout[57] ,\inst_twentynm_pma|w_pma_rx_deser_dout[56] ,\inst_twentynm_pma|w_pma_rx_deser_dout[55] ,\inst_twentynm_pma|w_pma_rx_deser_dout[54] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[53] ,\inst_twentynm_pma|w_pma_rx_deser_dout[52] ,\inst_twentynm_pma|w_pma_rx_deser_dout[51] ,\inst_twentynm_pma|w_pma_rx_deser_dout[50] ,\inst_twentynm_pma|w_pma_rx_deser_dout[49] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[48] ,\inst_twentynm_pma|w_pma_rx_deser_dout[47] ,\inst_twentynm_pma|w_pma_rx_deser_dout[46] ,\inst_twentynm_pma|w_pma_rx_deser_dout[45] ,\inst_twentynm_pma|w_pma_rx_deser_dout[44] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[43] ,\inst_twentynm_pma|w_pma_rx_deser_dout[42] ,\inst_twentynm_pma|w_pma_rx_deser_dout[41] ,\inst_twentynm_pma|w_pma_rx_deser_dout[40] ,\inst_twentynm_pma|w_pma_rx_deser_dout[39] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[38] ,\inst_twentynm_pma|w_pma_rx_deser_dout[37] ,\inst_twentynm_pma|w_pma_rx_deser_dout[36] ,\inst_twentynm_pma|w_pma_rx_deser_dout[35] ,\inst_twentynm_pma|w_pma_rx_deser_dout[34] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[33] ,\inst_twentynm_pma|w_pma_rx_deser_dout[32] ,\inst_twentynm_pma|w_pma_rx_deser_dout[31] ,\inst_twentynm_pma|w_pma_rx_deser_dout[30] ,\inst_twentynm_pma|w_pma_rx_deser_dout[29] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[28] ,\inst_twentynm_pma|w_pma_rx_deser_dout[27] ,\inst_twentynm_pma|w_pma_rx_deser_dout[26] ,\inst_twentynm_pma|w_pma_rx_deser_dout[25] ,\inst_twentynm_pma|w_pma_rx_deser_dout[24] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[23] ,\inst_twentynm_pma|w_pma_rx_deser_dout[22] ,\inst_twentynm_pma|w_pma_rx_deser_dout[21] ,\inst_twentynm_pma|w_pma_rx_deser_dout[20] ,\inst_twentynm_pma|w_pma_rx_deser_dout[19] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[18] ,\inst_twentynm_pma|w_pma_rx_deser_dout[17] ,\inst_twentynm_pma|w_pma_rx_deser_dout[16] ,\inst_twentynm_pma|w_pma_rx_deser_dout[15] ,\inst_twentynm_pma|w_pma_rx_deser_dout[14] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[13] ,\inst_twentynm_pma|w_pma_rx_deser_dout[12] ,\inst_twentynm_pma|w_pma_rx_deser_dout[11] ,\inst_twentynm_pma|w_pma_rx_deser_dout[10] ,\inst_twentynm_pma|w_pma_rx_deser_dout[9] ,\inst_twentynm_pma|w_pma_rx_deser_dout[8] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[7] ,\inst_twentynm_pma|w_pma_rx_deser_dout[6] ,\inst_twentynm_pma|w_pma_rx_deser_dout[5] ,\inst_twentynm_pma|w_pma_rx_deser_dout[4] ,\inst_twentynm_pma|w_pma_rx_deser_dout[3] ,\inst_twentynm_pma|w_pma_rx_deser_dout[2] ,
\inst_twentynm_pma|w_pma_rx_deser_dout[1] ,\inst_twentynm_pma|w_pma_rx_deser_dout[0] }),
	.out_blockselect_pma_rx_buf(\inst_twentynm_pma|w_pma_rx_buf_blockselect ),
	.out_avmmreaddata_pma_rx_buf({\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_buf_avmmreaddata[0] }),
	.out_blockselect_pma_rx_sd(\inst_twentynm_pma|w_pma_rx_sd_blockselect ),
	.out_sd(\inst_twentynm_pma|w_pma_rx_sd_sd ),
	.out_avmmreaddata_pma_rx_sd({\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_sd_avmmreaddata[0] }),
	.out_blockselect_pma_rx_odi(\inst_twentynm_pma|w_pma_rx_odi_blockselect ),
	.out_avmmreaddata_pma_rx_odi({\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_odi_avmmreaddata[0] }),
	.out_blockselect_pma_rx_dfe(\inst_twentynm_pma|w_pma_rx_dfe_blockselect ),
	.out_avmmreaddata_pma_rx_dfe({\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_rx_dfe_avmmreaddata[0] }),
	.out_blockselect_cdr_pll(\inst_twentynm_pma|w_cdr_pll_blockselect ),
	.out_clklow(\inst_twentynm_pma|w_cdr_pll_clklow ),
	.out_fref(\inst_twentynm_pma|w_cdr_pll_fref ),
	.out_pfdmode_lock(\inst_twentynm_pma|w_cdr_pll_pfdmode_lock ),
	.out_rxpll_lock(\inst_twentynm_pma|w_cdr_pll_rxpll_lock ),
	.out_avmmreaddata_cdr_pll({\inst_twentynm_pma|w_cdr_pll_avmmreaddata[7] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[6] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[5] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[4] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[3] ,
\inst_twentynm_pma|w_cdr_pll_avmmreaddata[2] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[1] ,\inst_twentynm_pma|w_cdr_pll_avmmreaddata[0] }),
	.out_blockselect_pma_cdr_refclk(\inst_twentynm_pma|w_pma_cdr_refclk_blockselect ),
	.out_avmmreaddata_pma_cdr_refclk({\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[4] ,
\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[3] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_cdr_refclk_avmmreaddata[0] }),
	.out_blockselect_pma_adapt(\inst_twentynm_pma|w_pma_adapt_blockselect ),
	.out_avmmreaddata_pma_adapt({\inst_twentynm_pma|w_pma_adapt_avmmreaddata[7] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[6] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[5] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[4] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[3] ,
\inst_twentynm_pma|w_pma_adapt_avmmreaddata[2] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[1] ,\inst_twentynm_pma|w_pma_adapt_avmmreaddata[0] }),
	.in_early_eios(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_early_eios ),
	.in_ltd_b(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltd_b ),
	.in_ltr(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ltr ),
	.in_ppm_lock(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_ppm_lock ),
	.in_rs_lpbk_b(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rs_lpbk_b ),
	.in_rx_qpi_pulldn(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_rx_qpi_pullup ),
	.in_tx_bitslip(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bitslip ),
	.in_tx_bonding_rstb(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_bonding_rstb ),
	.in_tx_qpi_pulldn(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pulldn ),
	.in_tx_qpi_pullup(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_qpi_pullup ),
	.in_tx_det_rx(\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_tx_txdetectrx ),
	.in_i_coeff({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[17] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[16] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[15] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[14] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[13] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[12] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[11] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[10] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[9] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[8] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[7] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[6] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[5] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[4] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[3] ,
\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[2] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_current_coeff[0] }),
	.in_pcie_sw({\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[1] ,\inst_twentynm_pcs|w_hssi_common_pcs_pma_interface_pma_pcie_switch[0] }),
	.in_tx_elec_idle(\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_elec_idle ),
	.in_tx_pma_rstb(\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_txpma_rstb ),
	.in_tx_data({\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[63] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[62] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[61] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[60] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[59] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[58] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[57] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[56] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[55] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[54] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[53] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[52] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[51] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[50] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[49] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[48] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[47] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[46] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[45] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[44] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[43] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[42] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[41] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[40] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[39] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[38] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[37] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[36] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[35] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[34] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[33] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[32] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[31] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[30] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[29] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[28] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[27] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[26] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[25] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[24] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[23] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[22] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[21] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[20] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[19] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[18] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[17] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[16] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[15] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[14] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[13] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[12] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[11] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[10] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[9] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[8] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[7] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[6] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[5] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[4] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[3] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[2] ,\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[1] ,
\inst_twentynm_pcs|w_hssi_tx_pcs_pma_interface_pma_tx_pma_data[0] }),
	.in_rx_p(rx_serial_data_0),
	.in_clk_fpll_b(tx_serial_clk0_0),
	.in_ref_iqclk({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rx_cdr_refclk0}));

endmodule

module wr_arria10_e3p1_det_phy_twentynm_pcs_rev_20nm5 (
	out_blockselect_hssi_rx_pld_pcs_interface,
	out_pld_pcs_rx_clk_out,
	out_avmmreaddata_hssi_rx_pld_pcs_interface,
	out_pld_8g_wa_boundary,
	out_pld_rx_data,
	in_avmmclk,
	in_avmmread,
	in_avmmrstn,
	in_avmmwrite,
	in_avmmaddress,
	in_avmmwritedata,
	out_blockselect_hssi_common_pld_pcs_interface,
	out_pld_pma_pfdmode_lock,
	out_pld_pma_rxpll_lock,
	out_avmmreaddata_hssi_common_pld_pcs_interface,
	out_blockselect_hssi_tx_pld_pcs_interface,
	out_pld_pcs_tx_clk_out,
	out_avmmreaddata_hssi_tx_pld_pcs_interface,
	in_pma_rx_detect_valid,
	in_pma_rx_found,
	out_blockselect_hssi_10g_rx_pcs,
	out_avmmreaddata_hssi_10g_rx_pcs,
	out_blockselect_hssi_8g_rx_pcs,
	out_avmmreaddata_hssi_8g_rx_pcs,
	out_blockselect_hssi_pipe_gen1_2,
	out_avmmreaddata_hssi_pipe_gen1_2,
	out_blockselect_hssi_krfec_rx_pcs,
	out_avmmreaddata_hssi_krfec_rx_pcs,
	out_blockselect_hssi_rx_pcs_pma_interface,
	out_pma_rx_clkslip,
	out_pma_rxpma_rstb,
	out_avmmreaddata_hssi_rx_pcs_pma_interface,
	out_pma_eye_monitor,
	in_pma_tx_pma_clk,
	in_pma_tx_clkdiv_user,
	in_pma_pcie_sw_done,
	in_pma_rx_pma_clk,
	in_pma_rx_clkdiv_user,
	in_pma_rx_pma_data,
	in_pma_signal_det,
	in_pma_clklow,
	in_pma_fref,
	in_pma_pfdmode_lock,
	in_pma_rxpll_lock,
	out_blockselect_hssi_8g_tx_pcs,
	out_avmmreaddata_hssi_8g_tx_pcs,
	out_blockselect_hssi_10g_tx_pcs,
	out_avmmreaddata_hssi_10g_tx_pcs,
	out_blockselect_hssi_gen3_rx_pcs,
	out_avmmreaddata_hssi_gen3_rx_pcs,
	out_blockselect_hssi_pipe_gen3,
	out_avmmreaddata_hssi_pipe_gen3,
	out_blockselect_hssi_gen3_tx_pcs,
	out_avmmreaddata_hssi_gen3_tx_pcs,
	out_blockselect_hssi_krfec_tx_pcs,
	out_avmmreaddata_hssi_krfec_tx_pcs,
	out_blockselect_hssi_fifo_rx_pcs,
	out_avmmreaddata_hssi_fifo_rx_pcs,
	out_blockselect_hssi_fifo_tx_pcs,
	out_avmmreaddata_hssi_fifo_tx_pcs,
	out_blockselect_hssi_common_pcs_pma_interface,
	out_pma_early_eios,
	out_pma_ltd_b,
	out_pma_ltr,
	out_pma_ppm_lock,
	out_pma_rs_lpbk_b,
	out_pma_rx_qpi_pullup,
	out_pma_tx_bitslip,
	out_pma_tx_bonding_rstb,
	out_pma_tx_qpi_pulldn,
	out_pma_tx_qpi_pullup,
	out_pma_tx_txdetectrx,
	out_avmmreaddata_hssi_common_pcs_pma_interface,
	out_pma_current_coeff,
	out_pma_pcie_switch,
	out_blockselect_hssi_tx_pcs_pma_interface,
	out_pma_tx_elec_idle,
	out_pma_txpma_rstb,
	out_avmmreaddata_hssi_tx_pcs_pma_interface,
	out_pma_tx_pma_data,
	in_pld_pma_txpma_rstb,
	in_pld_pma_rxpma_rstb,
	in_pld_10g_krfec_rx_pld_rst_n,
	in_pld_8g_g3_rx_pld_rst_n,
	in_pld_pmaif_rx_pld_rst_n,
	in_pld_8g_encdt,
	in_pld_rx_clk,
	in_pld_pma_rs_lpbk_b,
	in_pld_10g_krfec_tx_pld_rst_n,
	in_pld_8g_g3_tx_pld_rst_n,
	in_pld_pmaif_tx_pld_rst_n,
	in_pld_tx_clk,
	in_pld_tx_data)/* synthesis synthesis_greybox=1 */;
output 	out_blockselect_hssi_rx_pld_pcs_interface;
output 	out_pld_pcs_rx_clk_out;
output 	[7:0] out_avmmreaddata_hssi_rx_pld_pcs_interface;
output 	[4:0] out_pld_8g_wa_boundary;
output 	[127:0] out_pld_rx_data;
input 	in_avmmclk;
input 	in_avmmread;
input 	in_avmmrstn;
input 	in_avmmwrite;
input 	[8:0] in_avmmaddress;
input 	[7:0] in_avmmwritedata;
output 	out_blockselect_hssi_common_pld_pcs_interface;
output 	out_pld_pma_pfdmode_lock;
output 	out_pld_pma_rxpll_lock;
output 	[7:0] out_avmmreaddata_hssi_common_pld_pcs_interface;
output 	out_blockselect_hssi_tx_pld_pcs_interface;
output 	out_pld_pcs_tx_clk_out;
output 	[7:0] out_avmmreaddata_hssi_tx_pld_pcs_interface;
input 	in_pma_rx_detect_valid;
input 	in_pma_rx_found;
output 	out_blockselect_hssi_10g_rx_pcs;
output 	[7:0] out_avmmreaddata_hssi_10g_rx_pcs;
output 	out_blockselect_hssi_8g_rx_pcs;
output 	[7:0] out_avmmreaddata_hssi_8g_rx_pcs;
output 	out_blockselect_hssi_pipe_gen1_2;
output 	[7:0] out_avmmreaddata_hssi_pipe_gen1_2;
output 	out_blockselect_hssi_krfec_rx_pcs;
output 	[7:0] out_avmmreaddata_hssi_krfec_rx_pcs;
output 	out_blockselect_hssi_rx_pcs_pma_interface;
output 	out_pma_rx_clkslip;
output 	out_pma_rxpma_rstb;
output 	[7:0] out_avmmreaddata_hssi_rx_pcs_pma_interface;
output 	[5:0] out_pma_eye_monitor;
input 	in_pma_tx_pma_clk;
input 	in_pma_tx_clkdiv_user;
input 	[1:0] in_pma_pcie_sw_done;
input 	in_pma_rx_pma_clk;
input 	in_pma_rx_clkdiv_user;
input 	[63:0] in_pma_rx_pma_data;
input 	in_pma_signal_det;
input 	in_pma_clklow;
input 	in_pma_fref;
input 	in_pma_pfdmode_lock;
input 	in_pma_rxpll_lock;
output 	out_blockselect_hssi_8g_tx_pcs;
output 	[7:0] out_avmmreaddata_hssi_8g_tx_pcs;
output 	out_blockselect_hssi_10g_tx_pcs;
output 	[7:0] out_avmmreaddata_hssi_10g_tx_pcs;
output 	out_blockselect_hssi_gen3_rx_pcs;
output 	[7:0] out_avmmreaddata_hssi_gen3_rx_pcs;
output 	out_blockselect_hssi_pipe_gen3;
output 	[7:0] out_avmmreaddata_hssi_pipe_gen3;
output 	out_blockselect_hssi_gen3_tx_pcs;
output 	[7:0] out_avmmreaddata_hssi_gen3_tx_pcs;
output 	out_blockselect_hssi_krfec_tx_pcs;
output 	[7:0] out_avmmreaddata_hssi_krfec_tx_pcs;
output 	out_blockselect_hssi_fifo_rx_pcs;
output 	[7:0] out_avmmreaddata_hssi_fifo_rx_pcs;
output 	out_blockselect_hssi_fifo_tx_pcs;
output 	[7:0] out_avmmreaddata_hssi_fifo_tx_pcs;
output 	out_blockselect_hssi_common_pcs_pma_interface;
output 	out_pma_early_eios;
output 	out_pma_ltd_b;
output 	out_pma_ltr;
output 	out_pma_ppm_lock;
output 	out_pma_rs_lpbk_b;
output 	out_pma_rx_qpi_pullup;
output 	out_pma_tx_bitslip;
output 	out_pma_tx_bonding_rstb;
output 	out_pma_tx_qpi_pulldn;
output 	out_pma_tx_qpi_pullup;
output 	out_pma_tx_txdetectrx;
output 	[7:0] out_avmmreaddata_hssi_common_pcs_pma_interface;
output 	[17:0] out_pma_current_coeff;
output 	[1:0] out_pma_pcie_switch;
output 	out_blockselect_hssi_tx_pcs_pma_interface;
output 	out_pma_tx_elec_idle;
output 	out_pma_txpma_rstb;
output 	[7:0] out_avmmreaddata_hssi_tx_pcs_pma_interface;
output 	[63:0] out_pma_tx_pma_data;
input 	in_pld_pma_txpma_rstb;
input 	in_pld_pma_rxpma_rstb;
input 	in_pld_10g_krfec_rx_pld_rst_n;
input 	in_pld_8g_g3_rx_pld_rst_n;
input 	in_pld_pmaif_rx_pld_rst_n;
input 	in_pld_8g_encdt;
input 	in_pld_rx_clk;
input 	in_pld_pma_rs_lpbk_b;
input 	in_pld_10g_krfec_tx_pld_rst_n;
input 	in_pld_8g_g3_tx_pld_rst_n;
input 	in_pld_pmaif_tx_pld_rst_n;
input 	in_pld_tx_clk;
input 	[127:0] in_pld_tx_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs~O_STA_RX_CLK2_BY2_1 ;
wire \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs~O_STA_TX_CLK2_BY2_1 ;
wire \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface~O_STA_PMA_HCLK_BY2 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT0 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT1 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT2 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT3 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT4 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT5 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT6 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT7 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT8 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT9 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT10 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT11 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT12 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT13 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT14 ;
wire \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT15 ;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr;
wire w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en;
wire w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx;
wire w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en;
wire w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters;
wire w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx;
wire w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip;
wire w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n;
wire w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr;
wire w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126] ;
wire \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127] ;
wire w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig;
wire w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig;
wire w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2;
wire w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig;
wire w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx;
wire w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig;
wire w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel;
wire w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in;
wire w_hssi_common_pld_pcs_interface_scan_mode_n;
wire \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0] ;
wire \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1] ;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n;
wire w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n;
wire w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb;
wire w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62] ;
wire \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63] ;
wire w_hssi_10g_rx_pcs_rx_align_val;
wire w_hssi_10g_rx_pcs_rx_blk_lock;
wire w_hssi_10g_rx_pcs_rx_clk_out;
wire w_hssi_10g_rx_pcs_rx_clk_out_pld_if;
wire w_hssi_10g_rx_pcs_rx_crc32_err;
wire w_hssi_10g_rx_pcs_rx_data_valid;
wire w_hssi_10g_rx_pcs_rx_dft_clk_out;
wire w_hssi_10g_rx_pcs_rx_empty;
wire w_hssi_10g_rx_pcs_rx_fec_clk;
wire w_hssi_10g_rx_pcs_rx_fifo_del;
wire w_hssi_10g_rx_pcs_rx_fifo_insert;
wire w_hssi_10g_rx_pcs_rx_fifo_wr_clk;
wire w_hssi_10g_rx_pcs_rx_fifo_wr_en;
wire w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n;
wire w_hssi_10g_rx_pcs_rx_frame_lock;
wire w_hssi_10g_rx_pcs_rx_hi_ber;
wire w_hssi_10g_rx_pcs_rx_master_clk;
wire w_hssi_10g_rx_pcs_rx_master_clk_rst_n;
wire w_hssi_10g_rx_pcs_rx_oflw_err;
wire w_hssi_10g_rx_pcs_rx_pempty;
wire w_hssi_10g_rx_pcs_rx_pfull;
wire w_hssi_10g_rx_pcs_rx_random_err;
wire w_hssi_10g_rx_pcs_rx_rx_frame;
wire \w_hssi_10g_rx_pcs_rx_control[0] ;
wire \w_hssi_10g_rx_pcs_rx_control[1] ;
wire \w_hssi_10g_rx_pcs_rx_control[2] ;
wire \w_hssi_10g_rx_pcs_rx_control[3] ;
wire \w_hssi_10g_rx_pcs_rx_control[4] ;
wire \w_hssi_10g_rx_pcs_rx_control[5] ;
wire \w_hssi_10g_rx_pcs_rx_control[6] ;
wire \w_hssi_10g_rx_pcs_rx_control[7] ;
wire \w_hssi_10g_rx_pcs_rx_control[8] ;
wire \w_hssi_10g_rx_pcs_rx_control[9] ;
wire \w_hssi_10g_rx_pcs_rx_control[10] ;
wire \w_hssi_10g_rx_pcs_rx_control[11] ;
wire \w_hssi_10g_rx_pcs_rx_control[12] ;
wire \w_hssi_10g_rx_pcs_rx_control[13] ;
wire \w_hssi_10g_rx_pcs_rx_control[14] ;
wire \w_hssi_10g_rx_pcs_rx_control[15] ;
wire \w_hssi_10g_rx_pcs_rx_control[16] ;
wire \w_hssi_10g_rx_pcs_rx_control[17] ;
wire \w_hssi_10g_rx_pcs_rx_control[18] ;
wire \w_hssi_10g_rx_pcs_rx_control[19] ;
wire \w_hssi_10g_rx_pcs_rx_data[0] ;
wire \w_hssi_10g_rx_pcs_rx_data[1] ;
wire \w_hssi_10g_rx_pcs_rx_data[2] ;
wire \w_hssi_10g_rx_pcs_rx_data[3] ;
wire \w_hssi_10g_rx_pcs_rx_data[4] ;
wire \w_hssi_10g_rx_pcs_rx_data[5] ;
wire \w_hssi_10g_rx_pcs_rx_data[6] ;
wire \w_hssi_10g_rx_pcs_rx_data[7] ;
wire \w_hssi_10g_rx_pcs_rx_data[8] ;
wire \w_hssi_10g_rx_pcs_rx_data[9] ;
wire \w_hssi_10g_rx_pcs_rx_data[10] ;
wire \w_hssi_10g_rx_pcs_rx_data[11] ;
wire \w_hssi_10g_rx_pcs_rx_data[12] ;
wire \w_hssi_10g_rx_pcs_rx_data[13] ;
wire \w_hssi_10g_rx_pcs_rx_data[14] ;
wire \w_hssi_10g_rx_pcs_rx_data[15] ;
wire \w_hssi_10g_rx_pcs_rx_data[16] ;
wire \w_hssi_10g_rx_pcs_rx_data[17] ;
wire \w_hssi_10g_rx_pcs_rx_data[18] ;
wire \w_hssi_10g_rx_pcs_rx_data[19] ;
wire \w_hssi_10g_rx_pcs_rx_data[20] ;
wire \w_hssi_10g_rx_pcs_rx_data[21] ;
wire \w_hssi_10g_rx_pcs_rx_data[22] ;
wire \w_hssi_10g_rx_pcs_rx_data[23] ;
wire \w_hssi_10g_rx_pcs_rx_data[24] ;
wire \w_hssi_10g_rx_pcs_rx_data[25] ;
wire \w_hssi_10g_rx_pcs_rx_data[26] ;
wire \w_hssi_10g_rx_pcs_rx_data[27] ;
wire \w_hssi_10g_rx_pcs_rx_data[28] ;
wire \w_hssi_10g_rx_pcs_rx_data[29] ;
wire \w_hssi_10g_rx_pcs_rx_data[30] ;
wire \w_hssi_10g_rx_pcs_rx_data[31] ;
wire \w_hssi_10g_rx_pcs_rx_data[32] ;
wire \w_hssi_10g_rx_pcs_rx_data[33] ;
wire \w_hssi_10g_rx_pcs_rx_data[34] ;
wire \w_hssi_10g_rx_pcs_rx_data[35] ;
wire \w_hssi_10g_rx_pcs_rx_data[36] ;
wire \w_hssi_10g_rx_pcs_rx_data[37] ;
wire \w_hssi_10g_rx_pcs_rx_data[38] ;
wire \w_hssi_10g_rx_pcs_rx_data[39] ;
wire \w_hssi_10g_rx_pcs_rx_data[40] ;
wire \w_hssi_10g_rx_pcs_rx_data[41] ;
wire \w_hssi_10g_rx_pcs_rx_data[42] ;
wire \w_hssi_10g_rx_pcs_rx_data[43] ;
wire \w_hssi_10g_rx_pcs_rx_data[44] ;
wire \w_hssi_10g_rx_pcs_rx_data[45] ;
wire \w_hssi_10g_rx_pcs_rx_data[46] ;
wire \w_hssi_10g_rx_pcs_rx_data[47] ;
wire \w_hssi_10g_rx_pcs_rx_data[48] ;
wire \w_hssi_10g_rx_pcs_rx_data[49] ;
wire \w_hssi_10g_rx_pcs_rx_data[50] ;
wire \w_hssi_10g_rx_pcs_rx_data[51] ;
wire \w_hssi_10g_rx_pcs_rx_data[52] ;
wire \w_hssi_10g_rx_pcs_rx_data[53] ;
wire \w_hssi_10g_rx_pcs_rx_data[54] ;
wire \w_hssi_10g_rx_pcs_rx_data[55] ;
wire \w_hssi_10g_rx_pcs_rx_data[56] ;
wire \w_hssi_10g_rx_pcs_rx_data[57] ;
wire \w_hssi_10g_rx_pcs_rx_data[58] ;
wire \w_hssi_10g_rx_pcs_rx_data[59] ;
wire \w_hssi_10g_rx_pcs_rx_data[60] ;
wire \w_hssi_10g_rx_pcs_rx_data[61] ;
wire \w_hssi_10g_rx_pcs_rx_data[62] ;
wire \w_hssi_10g_rx_pcs_rx_data[63] ;
wire \w_hssi_10g_rx_pcs_rx_data[64] ;
wire \w_hssi_10g_rx_pcs_rx_data[65] ;
wire \w_hssi_10g_rx_pcs_rx_data[66] ;
wire \w_hssi_10g_rx_pcs_rx_data[67] ;
wire \w_hssi_10g_rx_pcs_rx_data[68] ;
wire \w_hssi_10g_rx_pcs_rx_data[69] ;
wire \w_hssi_10g_rx_pcs_rx_data[70] ;
wire \w_hssi_10g_rx_pcs_rx_data[71] ;
wire \w_hssi_10g_rx_pcs_rx_data[72] ;
wire \w_hssi_10g_rx_pcs_rx_data[73] ;
wire \w_hssi_10g_rx_pcs_rx_data[74] ;
wire \w_hssi_10g_rx_pcs_rx_data[75] ;
wire \w_hssi_10g_rx_pcs_rx_data[76] ;
wire \w_hssi_10g_rx_pcs_rx_data[77] ;
wire \w_hssi_10g_rx_pcs_rx_data[78] ;
wire \w_hssi_10g_rx_pcs_rx_data[79] ;
wire \w_hssi_10g_rx_pcs_rx_data[80] ;
wire \w_hssi_10g_rx_pcs_rx_data[81] ;
wire \w_hssi_10g_rx_pcs_rx_data[82] ;
wire \w_hssi_10g_rx_pcs_rx_data[83] ;
wire \w_hssi_10g_rx_pcs_rx_data[84] ;
wire \w_hssi_10g_rx_pcs_rx_data[85] ;
wire \w_hssi_10g_rx_pcs_rx_data[86] ;
wire \w_hssi_10g_rx_pcs_rx_data[87] ;
wire \w_hssi_10g_rx_pcs_rx_data[88] ;
wire \w_hssi_10g_rx_pcs_rx_data[89] ;
wire \w_hssi_10g_rx_pcs_rx_data[90] ;
wire \w_hssi_10g_rx_pcs_rx_data[91] ;
wire \w_hssi_10g_rx_pcs_rx_data[92] ;
wire \w_hssi_10g_rx_pcs_rx_data[93] ;
wire \w_hssi_10g_rx_pcs_rx_data[94] ;
wire \w_hssi_10g_rx_pcs_rx_data[95] ;
wire \w_hssi_10g_rx_pcs_rx_data[96] ;
wire \w_hssi_10g_rx_pcs_rx_data[97] ;
wire \w_hssi_10g_rx_pcs_rx_data[98] ;
wire \w_hssi_10g_rx_pcs_rx_data[99] ;
wire \w_hssi_10g_rx_pcs_rx_data[100] ;
wire \w_hssi_10g_rx_pcs_rx_data[101] ;
wire \w_hssi_10g_rx_pcs_rx_data[102] ;
wire \w_hssi_10g_rx_pcs_rx_data[103] ;
wire \w_hssi_10g_rx_pcs_rx_data[104] ;
wire \w_hssi_10g_rx_pcs_rx_data[105] ;
wire \w_hssi_10g_rx_pcs_rx_data[106] ;
wire \w_hssi_10g_rx_pcs_rx_data[107] ;
wire \w_hssi_10g_rx_pcs_rx_data[108] ;
wire \w_hssi_10g_rx_pcs_rx_data[109] ;
wire \w_hssi_10g_rx_pcs_rx_data[110] ;
wire \w_hssi_10g_rx_pcs_rx_data[111] ;
wire \w_hssi_10g_rx_pcs_rx_data[112] ;
wire \w_hssi_10g_rx_pcs_rx_data[113] ;
wire \w_hssi_10g_rx_pcs_rx_data[114] ;
wire \w_hssi_10g_rx_pcs_rx_data[115] ;
wire \w_hssi_10g_rx_pcs_rx_data[116] ;
wire \w_hssi_10g_rx_pcs_rx_data[117] ;
wire \w_hssi_10g_rx_pcs_rx_data[118] ;
wire \w_hssi_10g_rx_pcs_rx_data[119] ;
wire \w_hssi_10g_rx_pcs_rx_data[120] ;
wire \w_hssi_10g_rx_pcs_rx_data[121] ;
wire \w_hssi_10g_rx_pcs_rx_data[122] ;
wire \w_hssi_10g_rx_pcs_rx_data[123] ;
wire \w_hssi_10g_rx_pcs_rx_data[124] ;
wire \w_hssi_10g_rx_pcs_rx_data[125] ;
wire \w_hssi_10g_rx_pcs_rx_data[126] ;
wire \w_hssi_10g_rx_pcs_rx_data[127] ;
wire \w_hssi_10g_rx_pcs_rx_diag_status[0] ;
wire \w_hssi_10g_rx_pcs_rx_diag_status[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_num[0] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_num[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_num[2] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_num[3] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_num[4] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[0] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[2] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[3] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[4] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[5] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[6] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[7] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[8] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[9] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[10] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[11] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[12] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[13] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[14] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[15] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[16] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[17] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[18] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[19] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[20] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[21] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[22] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[23] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[24] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[25] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[26] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[27] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[28] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[29] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[30] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[31] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[32] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[33] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[34] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[35] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[36] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[37] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[38] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[39] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[40] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[41] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[42] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[43] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[44] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[45] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[46] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[47] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[48] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[49] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[50] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[51] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[52] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[53] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[54] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[55] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[56] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[57] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[58] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[59] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[60] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[61] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[62] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[63] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[64] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[65] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[66] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[67] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[68] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[69] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[70] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[71] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[72] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_data[73] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30] ;
wire \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31] ;
wire w_hssi_8g_rx_pcs_clock_to_pld;
wire w_hssi_8g_rx_pcs_dis_pc_byte;
wire w_hssi_8g_rx_pcs_eidle_detected;
wire w_hssi_8g_rx_pcs_g3_rx_pma_rstn;
wire w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn;
wire w_hssi_8g_rx_pcs_gen2ngen1;
wire w_hssi_8g_rx_pcs_pc_fifo_empty;
wire w_hssi_8g_rx_pcs_pcfifofull;
wire w_hssi_8g_rx_pcs_phystatus;
wire w_hssi_8g_rx_pcs_reset_pc_ptrs;
wire w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe;
wire w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe;
wire w_hssi_8g_rx_pcs_rm_fifo_empty;
wire w_hssi_8g_rx_pcs_rm_fifo_full;
wire w_hssi_8g_rx_pcs_rx_clk_out_pld_if;
wire w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if;
wire w_hssi_8g_rx_pcs_rx_clkslip;
wire w_hssi_8g_rx_pcs_rx_pipe_clk;
wire w_hssi_8g_rx_pcs_rx_pipe_soft_reset;
wire w_hssi_8g_rx_pcs_rx_pma_clk_gen3;
wire w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3;
wire w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g;
wire w_hssi_8g_rx_pcs_rxvalid;
wire w_hssi_8g_rx_pcs_signal_detect_out;
wire w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk;
wire w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk;
wire w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk;
wire w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk;
wire w_hssi_8g_rx_pcs_wr_en_rx_phfifo;
wire w_hssi_8g_rx_pcs_wr_en_rx_rmfifo;
wire w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo;
wire w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo;
wire \w_hssi_8g_rx_pcs_a1a2k1k2flag[0] ;
wire \w_hssi_8g_rx_pcs_a1a2k1k2flag[1] ;
wire \w_hssi_8g_rx_pcs_a1a2k1k2flag[2] ;
wire \w_hssi_8g_rx_pcs_a1a2k1k2flag[3] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[0] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[1] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[2] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[3] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[4] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[5] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[6] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[7] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[8] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[9] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[10] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[11] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[12] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[13] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[14] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[15] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[16] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[17] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[18] ;
wire \w_hssi_8g_rx_pcs_chnl_test_bus_out[19] ;
wire \w_hssi_8g_rx_pcs_dataout[0] ;
wire \w_hssi_8g_rx_pcs_dataout[1] ;
wire \w_hssi_8g_rx_pcs_dataout[2] ;
wire \w_hssi_8g_rx_pcs_dataout[3] ;
wire \w_hssi_8g_rx_pcs_dataout[4] ;
wire \w_hssi_8g_rx_pcs_dataout[5] ;
wire \w_hssi_8g_rx_pcs_dataout[6] ;
wire \w_hssi_8g_rx_pcs_dataout[7] ;
wire \w_hssi_8g_rx_pcs_dataout[8] ;
wire \w_hssi_8g_rx_pcs_dataout[9] ;
wire \w_hssi_8g_rx_pcs_dataout[10] ;
wire \w_hssi_8g_rx_pcs_dataout[11] ;
wire \w_hssi_8g_rx_pcs_dataout[12] ;
wire \w_hssi_8g_rx_pcs_dataout[13] ;
wire \w_hssi_8g_rx_pcs_dataout[14] ;
wire \w_hssi_8g_rx_pcs_dataout[15] ;
wire \w_hssi_8g_rx_pcs_dataout[16] ;
wire \w_hssi_8g_rx_pcs_dataout[17] ;
wire \w_hssi_8g_rx_pcs_dataout[18] ;
wire \w_hssi_8g_rx_pcs_dataout[19] ;
wire \w_hssi_8g_rx_pcs_dataout[20] ;
wire \w_hssi_8g_rx_pcs_dataout[21] ;
wire \w_hssi_8g_rx_pcs_dataout[22] ;
wire \w_hssi_8g_rx_pcs_dataout[23] ;
wire \w_hssi_8g_rx_pcs_dataout[24] ;
wire \w_hssi_8g_rx_pcs_dataout[25] ;
wire \w_hssi_8g_rx_pcs_dataout[26] ;
wire \w_hssi_8g_rx_pcs_dataout[27] ;
wire \w_hssi_8g_rx_pcs_dataout[28] ;
wire \w_hssi_8g_rx_pcs_dataout[29] ;
wire \w_hssi_8g_rx_pcs_dataout[30] ;
wire \w_hssi_8g_rx_pcs_dataout[31] ;
wire \w_hssi_8g_rx_pcs_dataout[32] ;
wire \w_hssi_8g_rx_pcs_dataout[33] ;
wire \w_hssi_8g_rx_pcs_dataout[34] ;
wire \w_hssi_8g_rx_pcs_dataout[35] ;
wire \w_hssi_8g_rx_pcs_dataout[36] ;
wire \w_hssi_8g_rx_pcs_dataout[37] ;
wire \w_hssi_8g_rx_pcs_dataout[38] ;
wire \w_hssi_8g_rx_pcs_dataout[39] ;
wire \w_hssi_8g_rx_pcs_dataout[40] ;
wire \w_hssi_8g_rx_pcs_dataout[41] ;
wire \w_hssi_8g_rx_pcs_dataout[42] ;
wire \w_hssi_8g_rx_pcs_dataout[43] ;
wire \w_hssi_8g_rx_pcs_dataout[44] ;
wire \w_hssi_8g_rx_pcs_dataout[45] ;
wire \w_hssi_8g_rx_pcs_dataout[46] ;
wire \w_hssi_8g_rx_pcs_dataout[47] ;
wire \w_hssi_8g_rx_pcs_dataout[48] ;
wire \w_hssi_8g_rx_pcs_dataout[49] ;
wire \w_hssi_8g_rx_pcs_dataout[50] ;
wire \w_hssi_8g_rx_pcs_dataout[51] ;
wire \w_hssi_8g_rx_pcs_dataout[52] ;
wire \w_hssi_8g_rx_pcs_dataout[53] ;
wire \w_hssi_8g_rx_pcs_dataout[54] ;
wire \w_hssi_8g_rx_pcs_dataout[55] ;
wire \w_hssi_8g_rx_pcs_dataout[56] ;
wire \w_hssi_8g_rx_pcs_dataout[57] ;
wire \w_hssi_8g_rx_pcs_dataout[58] ;
wire \w_hssi_8g_rx_pcs_dataout[59] ;
wire \w_hssi_8g_rx_pcs_dataout[60] ;
wire \w_hssi_8g_rx_pcs_dataout[61] ;
wire \w_hssi_8g_rx_pcs_dataout[62] ;
wire \w_hssi_8g_rx_pcs_dataout[63] ;
wire \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0] ;
wire \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1] ;
wire \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[0] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[1] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[2] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[3] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[4] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[5] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[6] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[7] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[8] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[9] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[10] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[11] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[12] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[13] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[14] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[15] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[16] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[17] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[18] ;
wire \w_hssi_8g_rx_pcs_parallel_rev_loopback[19] ;
wire \w_hssi_8g_rx_pcs_pipe_data[0] ;
wire \w_hssi_8g_rx_pcs_pipe_data[1] ;
wire \w_hssi_8g_rx_pcs_pipe_data[2] ;
wire \w_hssi_8g_rx_pcs_pipe_data[3] ;
wire \w_hssi_8g_rx_pcs_pipe_data[4] ;
wire \w_hssi_8g_rx_pcs_pipe_data[5] ;
wire \w_hssi_8g_rx_pcs_pipe_data[6] ;
wire \w_hssi_8g_rx_pcs_pipe_data[7] ;
wire \w_hssi_8g_rx_pcs_pipe_data[8] ;
wire \w_hssi_8g_rx_pcs_pipe_data[9] ;
wire \w_hssi_8g_rx_pcs_pipe_data[10] ;
wire \w_hssi_8g_rx_pcs_pipe_data[11] ;
wire \w_hssi_8g_rx_pcs_pipe_data[12] ;
wire \w_hssi_8g_rx_pcs_pipe_data[13] ;
wire \w_hssi_8g_rx_pcs_pipe_data[14] ;
wire \w_hssi_8g_rx_pcs_pipe_data[15] ;
wire \w_hssi_8g_rx_pcs_pipe_data[16] ;
wire \w_hssi_8g_rx_pcs_pipe_data[17] ;
wire \w_hssi_8g_rx_pcs_pipe_data[18] ;
wire \w_hssi_8g_rx_pcs_pipe_data[19] ;
wire \w_hssi_8g_rx_pcs_pipe_data[20] ;
wire \w_hssi_8g_rx_pcs_pipe_data[21] ;
wire \w_hssi_8g_rx_pcs_pipe_data[22] ;
wire \w_hssi_8g_rx_pcs_pipe_data[23] ;
wire \w_hssi_8g_rx_pcs_pipe_data[24] ;
wire \w_hssi_8g_rx_pcs_pipe_data[25] ;
wire \w_hssi_8g_rx_pcs_pipe_data[26] ;
wire \w_hssi_8g_rx_pcs_pipe_data[27] ;
wire \w_hssi_8g_rx_pcs_pipe_data[28] ;
wire \w_hssi_8g_rx_pcs_pipe_data[29] ;
wire \w_hssi_8g_rx_pcs_pipe_data[30] ;
wire \w_hssi_8g_rx_pcs_pipe_data[31] ;
wire \w_hssi_8g_rx_pcs_pipe_data[32] ;
wire \w_hssi_8g_rx_pcs_pipe_data[33] ;
wire \w_hssi_8g_rx_pcs_pipe_data[34] ;
wire \w_hssi_8g_rx_pcs_pipe_data[35] ;
wire \w_hssi_8g_rx_pcs_pipe_data[36] ;
wire \w_hssi_8g_rx_pcs_pipe_data[37] ;
wire \w_hssi_8g_rx_pcs_pipe_data[38] ;
wire \w_hssi_8g_rx_pcs_pipe_data[39] ;
wire \w_hssi_8g_rx_pcs_pipe_data[40] ;
wire \w_hssi_8g_rx_pcs_pipe_data[41] ;
wire \w_hssi_8g_rx_pcs_pipe_data[42] ;
wire \w_hssi_8g_rx_pcs_pipe_data[43] ;
wire \w_hssi_8g_rx_pcs_pipe_data[44] ;
wire \w_hssi_8g_rx_pcs_pipe_data[45] ;
wire \w_hssi_8g_rx_pcs_pipe_data[46] ;
wire \w_hssi_8g_rx_pcs_pipe_data[47] ;
wire \w_hssi_8g_rx_pcs_pipe_data[48] ;
wire \w_hssi_8g_rx_pcs_pipe_data[49] ;
wire \w_hssi_8g_rx_pcs_pipe_data[50] ;
wire \w_hssi_8g_rx_pcs_pipe_data[51] ;
wire \w_hssi_8g_rx_pcs_pipe_data[52] ;
wire \w_hssi_8g_rx_pcs_pipe_data[53] ;
wire \w_hssi_8g_rx_pcs_pipe_data[54] ;
wire \w_hssi_8g_rx_pcs_pipe_data[55] ;
wire \w_hssi_8g_rx_pcs_pipe_data[56] ;
wire \w_hssi_8g_rx_pcs_pipe_data[57] ;
wire \w_hssi_8g_rx_pcs_pipe_data[58] ;
wire \w_hssi_8g_rx_pcs_pipe_data[59] ;
wire \w_hssi_8g_rx_pcs_pipe_data[60] ;
wire \w_hssi_8g_rx_pcs_pipe_data[61] ;
wire \w_hssi_8g_rx_pcs_pipe_data[62] ;
wire \w_hssi_8g_rx_pcs_pipe_data[63] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18] ;
wire \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18] ;
wire \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6] ;
wire \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7] ;
wire \w_hssi_8g_rx_pcs_rx_blk_start[0] ;
wire \w_hssi_8g_rx_pcs_rx_blk_start[1] ;
wire \w_hssi_8g_rx_pcs_rx_blk_start[2] ;
wire \w_hssi_8g_rx_pcs_rx_blk_start[3] ;
wire \w_hssi_8g_rx_pcs_rx_data_valid[0] ;
wire \w_hssi_8g_rx_pcs_rx_data_valid[1] ;
wire \w_hssi_8g_rx_pcs_rx_data_valid[2] ;
wire \w_hssi_8g_rx_pcs_rx_data_valid[3] ;
wire \w_hssi_8g_rx_pcs_rx_sync_hdr[0] ;
wire \w_hssi_8g_rx_pcs_rx_sync_hdr[1] ;
wire \w_hssi_8g_rx_pcs_rxstatus[0] ;
wire \w_hssi_8g_rx_pcs_rxstatus[1] ;
wire \w_hssi_8g_rx_pcs_rxstatus[2] ;
wire \w_hssi_8g_rx_pcs_word_align_boundary[0] ;
wire \w_hssi_8g_rx_pcs_word_align_boundary[1] ;
wire \w_hssi_8g_rx_pcs_word_align_boundary[2] ;
wire \w_hssi_8g_rx_pcs_word_align_boundary[3] ;
wire \w_hssi_8g_rx_pcs_word_align_boundary[4] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30] ;
wire \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18] ;
wire \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19] ;
wire w_hssi_pipe_gen1_2_phystatus;
wire w_hssi_pipe_gen1_2_polarity_inversion_rx;
wire w_hssi_pipe_gen1_2_rev_loopbk;
wire w_hssi_pipe_gen1_2_rxelecidle;
wire w_hssi_pipe_gen1_2_rxelectricalidle_out;
wire w_hssi_pipe_gen1_2_rxvalid;
wire w_hssi_pipe_gen1_2_tx_elec_idle_out;
wire w_hssi_pipe_gen1_2_txdetectrx;
wire \w_hssi_pipe_gen1_2_current_coeff[0] ;
wire \w_hssi_pipe_gen1_2_current_coeff[1] ;
wire \w_hssi_pipe_gen1_2_current_coeff[2] ;
wire \w_hssi_pipe_gen1_2_current_coeff[3] ;
wire \w_hssi_pipe_gen1_2_current_coeff[4] ;
wire \w_hssi_pipe_gen1_2_current_coeff[5] ;
wire \w_hssi_pipe_gen1_2_current_coeff[6] ;
wire \w_hssi_pipe_gen1_2_current_coeff[7] ;
wire \w_hssi_pipe_gen1_2_current_coeff[8] ;
wire \w_hssi_pipe_gen1_2_current_coeff[9] ;
wire \w_hssi_pipe_gen1_2_current_coeff[10] ;
wire \w_hssi_pipe_gen1_2_current_coeff[11] ;
wire \w_hssi_pipe_gen1_2_current_coeff[12] ;
wire \w_hssi_pipe_gen1_2_current_coeff[13] ;
wire \w_hssi_pipe_gen1_2_current_coeff[14] ;
wire \w_hssi_pipe_gen1_2_current_coeff[15] ;
wire \w_hssi_pipe_gen1_2_current_coeff[16] ;
wire \w_hssi_pipe_gen1_2_current_coeff[17] ;
wire \w_hssi_pipe_gen1_2_rxstatus[0] ;
wire \w_hssi_pipe_gen1_2_rxstatus[1] ;
wire \w_hssi_pipe_gen1_2_rxstatus[2] ;
wire w_hssi_krfec_rx_pcs_rx_block_lock;
wire w_hssi_krfec_rx_pcs_rx_data_valid_out;
wire w_hssi_krfec_rx_pcs_rx_frame;
wire w_hssi_krfec_rx_pcs_rx_signal_ok_out;
wire \w_hssi_krfec_rx_pcs_rx_control_out[0] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[1] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[2] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[3] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[4] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[5] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[6] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[7] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[8] ;
wire \w_hssi_krfec_rx_pcs_rx_control_out[9] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[0] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[1] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[2] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[3] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[4] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[5] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[6] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[7] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[8] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[9] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[10] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[11] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[12] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[13] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[14] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[15] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[16] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[17] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[18] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[19] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[20] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[21] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[22] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[23] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[24] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[25] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[26] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[27] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[28] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[29] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[30] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[31] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[32] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[33] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[34] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[35] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[36] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[37] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[38] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[39] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[40] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[41] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[42] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[43] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[44] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[45] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[46] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[47] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[48] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[49] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[50] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[51] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[52] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[53] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[54] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[55] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[56] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[57] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[58] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[59] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[60] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[61] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[62] ;
wire \w_hssi_krfec_rx_pcs_rx_data_out[63] ;
wire \w_hssi_krfec_rx_pcs_rx_data_status[0] ;
wire \w_hssi_krfec_rx_pcs_rx_data_status[1] ;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock;
wire w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok;
wire w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62] ;
wire \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18] ;
wire \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18] ;
wire \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19] ;
wire w_hssi_8g_tx_pcs_clk_out;
wire w_hssi_8g_tx_pcs_clk_out_gen3;
wire w_hssi_8g_tx_pcs_dyn_clk_switch_n;
wire w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn;
wire w_hssi_8g_tx_pcs_g3_tx_pma_rstn;
wire w_hssi_8g_tx_pcs_ph_fifo_overflow;
wire w_hssi_8g_tx_pcs_ph_fifo_underflow;
wire w_hssi_8g_tx_pcs_phfifo_txdeemph;
wire w_hssi_8g_tx_pcs_phfifo_txswing;
wire w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out;
wire w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3;
wire w_hssi_8g_tx_pcs_pmaif_asn_rstn;
wire w_hssi_8g_tx_pcs_refclk_b;
wire w_hssi_8g_tx_pcs_refclk_b_reset;
wire w_hssi_8g_tx_pcs_rxpolarity_int;
wire w_hssi_8g_tx_pcs_soft_reset_wclk1_n;
wire w_hssi_8g_tx_pcs_sw_fifo_wr_clk;
wire w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif;
wire w_hssi_8g_tx_pcs_tx_clk_out_pld_if;
wire w_hssi_8g_tx_pcs_tx_clk_out_pmaif;
wire w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if;
wire w_hssi_8g_tx_pcs_tx_detect_rxloopback_int;
wire w_hssi_8g_tx_pcs_tx_pipe_clk;
wire w_hssi_8g_tx_pcs_tx_pipe_electidle;
wire w_hssi_8g_tx_pcs_tx_pipe_soft_reset;
wire w_hssi_8g_tx_pcs_txcompliance_out;
wire w_hssi_8g_tx_pcs_txelecidle_out;
wire w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk;
wire w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk;
wire w_hssi_8g_tx_pcs_wr_en_tx_phfifo;
wire w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo;
wire \w_hssi_8g_tx_pcs_dataout[0] ;
wire \w_hssi_8g_tx_pcs_dataout[1] ;
wire \w_hssi_8g_tx_pcs_dataout[2] ;
wire \w_hssi_8g_tx_pcs_dataout[3] ;
wire \w_hssi_8g_tx_pcs_dataout[4] ;
wire \w_hssi_8g_tx_pcs_dataout[5] ;
wire \w_hssi_8g_tx_pcs_dataout[6] ;
wire \w_hssi_8g_tx_pcs_dataout[7] ;
wire \w_hssi_8g_tx_pcs_dataout[8] ;
wire \w_hssi_8g_tx_pcs_dataout[9] ;
wire \w_hssi_8g_tx_pcs_dataout[10] ;
wire \w_hssi_8g_tx_pcs_dataout[11] ;
wire \w_hssi_8g_tx_pcs_dataout[12] ;
wire \w_hssi_8g_tx_pcs_dataout[13] ;
wire \w_hssi_8g_tx_pcs_dataout[14] ;
wire \w_hssi_8g_tx_pcs_dataout[15] ;
wire \w_hssi_8g_tx_pcs_dataout[16] ;
wire \w_hssi_8g_tx_pcs_dataout[17] ;
wire \w_hssi_8g_tx_pcs_dataout[18] ;
wire \w_hssi_8g_tx_pcs_dataout[19] ;
wire \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0] ;
wire \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1] ;
wire \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2] ;
wire \w_hssi_8g_tx_pcs_phfifo_txmargin[0] ;
wire \w_hssi_8g_tx_pcs_phfifo_txmargin[1] ;
wire \w_hssi_8g_tx_pcs_phfifo_txmargin[2] ;
wire \w_hssi_8g_tx_pcs_pipe_power_down_out[0] ;
wire \w_hssi_8g_tx_pcs_pipe_power_down_out[1] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6] ;
wire \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7] ;
wire \w_hssi_8g_tx_pcs_tx_blk_start_out[0] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18] ;
wire \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[0] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[1] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[2] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[3] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[4] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[5] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[6] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[7] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[8] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[9] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[10] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[11] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[12] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[13] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[14] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[15] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[16] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[17] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[18] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[19] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[20] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[21] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[22] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[23] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[24] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[25] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[26] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[27] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[28] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[29] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[30] ;
wire \w_hssi_8g_tx_pcs_tx_data_out[31] ;
wire \w_hssi_8g_tx_pcs_tx_data_valid_out[0] ;
wire \w_hssi_8g_tx_pcs_tx_datak_out[0] ;
wire \w_hssi_8g_tx_pcs_tx_datak_out[1] ;
wire \w_hssi_8g_tx_pcs_tx_datak_out[2] ;
wire \w_hssi_8g_tx_pcs_tx_datak_out[3] ;
wire \w_hssi_8g_tx_pcs_tx_div_sync[0] ;
wire \w_hssi_8g_tx_pcs_tx_div_sync[1] ;
wire \w_hssi_8g_tx_pcs_tx_sync_hdr_out[0] ;
wire \w_hssi_8g_tx_pcs_tx_sync_hdr_out[1] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[0] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[1] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[2] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[3] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[4] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[5] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[6] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[7] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[8] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[9] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[10] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[11] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[12] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[13] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[14] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[15] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[16] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[17] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[18] ;
wire \w_hssi_8g_tx_pcs_tx_testbus[19] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62] ;
wire \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6] ;
wire \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7] ;
wire w_hssi_10g_tx_pcs_tx_burst_en_exe;
wire w_hssi_10g_tx_pcs_tx_clk_out;
wire w_hssi_10g_tx_pcs_tx_clk_out_pld_if;
wire w_hssi_10g_tx_pcs_tx_clk_out_pma_if;
wire w_hssi_10g_tx_pcs_tx_data_valid_out_krfec;
wire w_hssi_10g_tx_pcs_tx_dft_clk_out;
wire w_hssi_10g_tx_pcs_tx_empty;
wire w_hssi_10g_tx_pcs_tx_fec_clk;
wire w_hssi_10g_tx_pcs_tx_fifo_wr_clk;
wire w_hssi_10g_tx_pcs_tx_fifo_wr_en;
wire w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n;
wire w_hssi_10g_tx_pcs_tx_frame;
wire w_hssi_10g_tx_pcs_tx_full;
wire w_hssi_10g_tx_pcs_tx_master_clk;
wire w_hssi_10g_tx_pcs_tx_master_clk_rst_n;
wire w_hssi_10g_tx_pcs_tx_pempty;
wire w_hssi_10g_tx_pcs_tx_pfull;
wire w_hssi_10g_tx_pcs_tx_wordslip_exe;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[0] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[1] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[2] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[3] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[4] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[5] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[6] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[7] ;
wire \w_hssi_10g_tx_pcs_tx_control_out_krfec[8] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[0] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[1] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[2] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[3] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[4] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[5] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[6] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[7] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[8] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[9] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[10] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[11] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[12] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[13] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[14] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[15] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[16] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[17] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[18] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[19] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[20] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[21] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[22] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[23] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[24] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[25] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[26] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[27] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[28] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[29] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[30] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[31] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[32] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[33] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[34] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[35] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[36] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[37] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[38] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[39] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[40] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[41] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[42] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[43] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[44] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[45] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[46] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[47] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[48] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[49] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[50] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[51] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[52] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[53] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[54] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[55] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[56] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[57] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[58] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[59] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[60] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[61] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[62] ;
wire \w_hssi_10g_tx_pcs_tx_data_out_krfec[63] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_num[0] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_num[1] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_num[2] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_num[3] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[0] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[1] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[2] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[3] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[4] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[5] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[6] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[7] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[8] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[9] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[10] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[11] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[12] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[13] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[14] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[15] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[16] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[17] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[18] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[19] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[20] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[21] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[22] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[23] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[24] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[25] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[26] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[27] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[28] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[29] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[30] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[31] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[32] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[33] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[34] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[35] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[36] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[37] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[38] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[39] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[40] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[41] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[42] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[43] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[44] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[45] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[46] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[47] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[48] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[49] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[50] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[51] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[52] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[53] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[54] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[55] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[56] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[57] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[58] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[59] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[60] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[61] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[62] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[63] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[64] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[65] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[66] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[67] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[68] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[69] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[70] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[71] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data[72] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14] ;
wire \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[0] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[1] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[2] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[3] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[4] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[5] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[6] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[7] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[8] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[9] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[10] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[11] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[12] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[13] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[14] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[15] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[16] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[17] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[18] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[19] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[20] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[21] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[22] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[23] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[24] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[25] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[26] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[27] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[28] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[29] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[30] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[31] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[32] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[33] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[34] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[35] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[36] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[37] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[38] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[39] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[40] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[41] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[42] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[43] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[44] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[45] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[46] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[47] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[48] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[49] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[50] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[51] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[52] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[53] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[54] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[55] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[56] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[57] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[58] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[59] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[60] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[61] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[62] ;
wire \w_hssi_10g_tx_pcs_tx_pma_data[63] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[0] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[1] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[2] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[3] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[4] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[5] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[6] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[7] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[8] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[9] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[10] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[11] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[12] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[13] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[14] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[15] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[16] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[17] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[18] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[19] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[20] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[21] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[22] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[23] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[24] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[25] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[26] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[27] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[28] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[29] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[30] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[31] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[32] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[33] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[34] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[35] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[36] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[37] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[38] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[39] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[40] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[41] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[42] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[43] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[44] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[45] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[46] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[47] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[48] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[49] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[50] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[51] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[52] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[53] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[54] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[55] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[56] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[57] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[58] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[59] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[60] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[61] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[62] ;
wire \w_hssi_10g_tx_pcs_tx_pma_gating_val[63] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[0] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[1] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[2] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[3] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[4] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[5] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[6] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[7] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[8] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[9] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[10] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[11] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[12] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[13] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[14] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[15] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[16] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[17] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[18] ;
wire \w_hssi_10g_tx_pcs_tx_test_data[19] ;
wire w_hssi_gen3_rx_pcs_blk_algnd_int;
wire w_hssi_gen3_rx_pcs_blk_start;
wire w_hssi_gen3_rx_pcs_clkcomp_delete_int;
wire w_hssi_gen3_rx_pcs_clkcomp_insert_int;
wire w_hssi_gen3_rx_pcs_clkcomp_overfl_int;
wire w_hssi_gen3_rx_pcs_clkcomp_undfl_int;
wire w_hssi_gen3_rx_pcs_data_valid;
wire w_hssi_gen3_rx_pcs_ei_det_int;
wire w_hssi_gen3_rx_pcs_ei_partial_det_int;
wire w_hssi_gen3_rx_pcs_err_decode_int;
wire w_hssi_gen3_rx_pcs_i_det_int;
wire w_hssi_gen3_rx_pcs_lpbk_blk_start;
wire w_hssi_gen3_rx_pcs_lpbk_data_valid;
wire w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk;
wire w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en;
wire w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n;
wire w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int;
wire \w_hssi_gen3_rx_pcs_data_out[0] ;
wire \w_hssi_gen3_rx_pcs_data_out[1] ;
wire \w_hssi_gen3_rx_pcs_data_out[2] ;
wire \w_hssi_gen3_rx_pcs_data_out[3] ;
wire \w_hssi_gen3_rx_pcs_data_out[4] ;
wire \w_hssi_gen3_rx_pcs_data_out[5] ;
wire \w_hssi_gen3_rx_pcs_data_out[6] ;
wire \w_hssi_gen3_rx_pcs_data_out[7] ;
wire \w_hssi_gen3_rx_pcs_data_out[8] ;
wire \w_hssi_gen3_rx_pcs_data_out[9] ;
wire \w_hssi_gen3_rx_pcs_data_out[10] ;
wire \w_hssi_gen3_rx_pcs_data_out[11] ;
wire \w_hssi_gen3_rx_pcs_data_out[12] ;
wire \w_hssi_gen3_rx_pcs_data_out[13] ;
wire \w_hssi_gen3_rx_pcs_data_out[14] ;
wire \w_hssi_gen3_rx_pcs_data_out[15] ;
wire \w_hssi_gen3_rx_pcs_data_out[16] ;
wire \w_hssi_gen3_rx_pcs_data_out[17] ;
wire \w_hssi_gen3_rx_pcs_data_out[18] ;
wire \w_hssi_gen3_rx_pcs_data_out[19] ;
wire \w_hssi_gen3_rx_pcs_data_out[20] ;
wire \w_hssi_gen3_rx_pcs_data_out[21] ;
wire \w_hssi_gen3_rx_pcs_data_out[22] ;
wire \w_hssi_gen3_rx_pcs_data_out[23] ;
wire \w_hssi_gen3_rx_pcs_data_out[24] ;
wire \w_hssi_gen3_rx_pcs_data_out[25] ;
wire \w_hssi_gen3_rx_pcs_data_out[26] ;
wire \w_hssi_gen3_rx_pcs_data_out[27] ;
wire \w_hssi_gen3_rx_pcs_data_out[28] ;
wire \w_hssi_gen3_rx_pcs_data_out[29] ;
wire \w_hssi_gen3_rx_pcs_data_out[30] ;
wire \w_hssi_gen3_rx_pcs_data_out[31] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[0] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[1] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[2] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[3] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[4] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[5] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[6] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[7] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[8] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[9] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[10] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[11] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[12] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[13] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[14] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[15] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[16] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[17] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[18] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[19] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[20] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[21] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[22] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[23] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[24] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[25] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[26] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[27] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[28] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[29] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[30] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[31] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[32] ;
wire \w_hssi_gen3_rx_pcs_lpbk_data[33] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14] ;
wire \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[0] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[1] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[2] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[3] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[4] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[5] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[6] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[7] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[8] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[9] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[10] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[11] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[12] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[13] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[14] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[15] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[16] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[17] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[18] ;
wire \w_hssi_gen3_rx_pcs_rx_test_out[19] ;
wire \w_hssi_gen3_rx_pcs_sync_hdr[0] ;
wire \w_hssi_gen3_rx_pcs_sync_hdr[1] ;
wire w_hssi_pipe_gen3_gen3_clk_sel;
wire w_hssi_pipe_gen3_pcs_rst;
wire w_hssi_pipe_gen3_phystatus;
wire w_hssi_pipe_gen3_pma_tx_elec_idle;
wire w_hssi_pipe_gen3_pma_txdetectrx;
wire w_hssi_pipe_gen3_rev_lpbk_8gpcs_out;
wire w_hssi_pipe_gen3_rev_lpbk_int;
wire w_hssi_pipe_gen3_rxelecidle;
wire w_hssi_pipe_gen3_rxpolarity_8gpcs_out;
wire w_hssi_pipe_gen3_rxpolarity_int;
wire w_hssi_pipe_gen3_rxvalid;
wire w_hssi_pipe_gen3_shutdown_clk;
wire w_hssi_pipe_gen3_tx_blk_start_int;
wire w_hssi_pipe_gen3_txdataskip_int;
wire \w_hssi_pipe_gen3_pma_current_coeff[0] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[1] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[2] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[3] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[4] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[5] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[6] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[7] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[8] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[9] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[10] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[11] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[12] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[13] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[14] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[15] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[16] ;
wire \w_hssi_pipe_gen3_pma_current_coeff[17] ;
wire \w_hssi_pipe_gen3_pma_current_rxpreset[0] ;
wire \w_hssi_pipe_gen3_pma_current_rxpreset[1] ;
wire \w_hssi_pipe_gen3_pma_current_rxpreset[2] ;
wire \w_hssi_pipe_gen3_rx_blk_start[0] ;
wire \w_hssi_pipe_gen3_rx_blk_start[1] ;
wire \w_hssi_pipe_gen3_rx_blk_start[2] ;
wire \w_hssi_pipe_gen3_rx_blk_start[3] ;
wire \w_hssi_pipe_gen3_rx_sync_hdr[0] ;
wire \w_hssi_pipe_gen3_rx_sync_hdr[1] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[0] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[1] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[2] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[3] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[4] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[5] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[6] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[7] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[8] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[9] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[10] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[11] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[12] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[13] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[14] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[15] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[16] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[17] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[18] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[19] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[20] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[21] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[22] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[23] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[24] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[25] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[26] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[27] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[28] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[29] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[30] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[31] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[32] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[33] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[34] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[35] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[36] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[37] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[38] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[39] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[40] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[41] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[42] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[43] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[44] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[45] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[46] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[47] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[48] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[49] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[50] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[51] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[52] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[53] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[54] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[55] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[56] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[57] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[58] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[59] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[60] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[61] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[62] ;
wire \w_hssi_pipe_gen3_rxd_8gpcs_out[63] ;
wire \w_hssi_pipe_gen3_rxdataskip[0] ;
wire \w_hssi_pipe_gen3_rxdataskip[1] ;
wire \w_hssi_pipe_gen3_rxdataskip[2] ;
wire \w_hssi_pipe_gen3_rxdataskip[3] ;
wire \w_hssi_pipe_gen3_rxstatus[0] ;
wire \w_hssi_pipe_gen3_rxstatus[1] ;
wire \w_hssi_pipe_gen3_rxstatus[2] ;
wire \w_hssi_pipe_gen3_test_out[0] ;
wire \w_hssi_pipe_gen3_test_out[1] ;
wire \w_hssi_pipe_gen3_test_out[2] ;
wire \w_hssi_pipe_gen3_test_out[3] ;
wire \w_hssi_pipe_gen3_test_out[4] ;
wire \w_hssi_pipe_gen3_test_out[5] ;
wire \w_hssi_pipe_gen3_test_out[6] ;
wire \w_hssi_pipe_gen3_test_out[7] ;
wire \w_hssi_pipe_gen3_test_out[8] ;
wire \w_hssi_pipe_gen3_test_out[9] ;
wire \w_hssi_pipe_gen3_test_out[10] ;
wire \w_hssi_pipe_gen3_test_out[11] ;
wire \w_hssi_pipe_gen3_test_out[12] ;
wire \w_hssi_pipe_gen3_test_out[13] ;
wire \w_hssi_pipe_gen3_test_out[14] ;
wire \w_hssi_pipe_gen3_test_out[15] ;
wire \w_hssi_pipe_gen3_test_out[16] ;
wire \w_hssi_pipe_gen3_test_out[17] ;
wire \w_hssi_pipe_gen3_test_out[18] ;
wire \w_hssi_pipe_gen3_test_out[19] ;
wire \w_hssi_pipe_gen3_tx_sync_hdr_int[0] ;
wire \w_hssi_pipe_gen3_tx_sync_hdr_int[1] ;
wire \w_hssi_pipe_gen3_txdata_int[0] ;
wire \w_hssi_pipe_gen3_txdata_int[1] ;
wire \w_hssi_pipe_gen3_txdata_int[2] ;
wire \w_hssi_pipe_gen3_txdata_int[3] ;
wire \w_hssi_pipe_gen3_txdata_int[4] ;
wire \w_hssi_pipe_gen3_txdata_int[5] ;
wire \w_hssi_pipe_gen3_txdata_int[6] ;
wire \w_hssi_pipe_gen3_txdata_int[7] ;
wire \w_hssi_pipe_gen3_txdata_int[8] ;
wire \w_hssi_pipe_gen3_txdata_int[9] ;
wire \w_hssi_pipe_gen3_txdata_int[10] ;
wire \w_hssi_pipe_gen3_txdata_int[11] ;
wire \w_hssi_pipe_gen3_txdata_int[12] ;
wire \w_hssi_pipe_gen3_txdata_int[13] ;
wire \w_hssi_pipe_gen3_txdata_int[14] ;
wire \w_hssi_pipe_gen3_txdata_int[15] ;
wire \w_hssi_pipe_gen3_txdata_int[16] ;
wire \w_hssi_pipe_gen3_txdata_int[17] ;
wire \w_hssi_pipe_gen3_txdata_int[18] ;
wire \w_hssi_pipe_gen3_txdata_int[19] ;
wire \w_hssi_pipe_gen3_txdata_int[20] ;
wire \w_hssi_pipe_gen3_txdata_int[21] ;
wire \w_hssi_pipe_gen3_txdata_int[22] ;
wire \w_hssi_pipe_gen3_txdata_int[23] ;
wire \w_hssi_pipe_gen3_txdata_int[24] ;
wire \w_hssi_pipe_gen3_txdata_int[25] ;
wire \w_hssi_pipe_gen3_txdata_int[26] ;
wire \w_hssi_pipe_gen3_txdata_int[27] ;
wire \w_hssi_pipe_gen3_txdata_int[28] ;
wire \w_hssi_pipe_gen3_txdata_int[29] ;
wire \w_hssi_pipe_gen3_txdata_int[30] ;
wire \w_hssi_pipe_gen3_txdata_int[31] ;
wire \w_hssi_pipe_gen3_txdatak_int[0] ;
wire \w_hssi_pipe_gen3_txdatak_int[1] ;
wire \w_hssi_pipe_gen3_txdatak_int[2] ;
wire \w_hssi_pipe_gen3_txdatak_int[3] ;
wire \w_hssi_gen3_tx_pcs_data_out[0] ;
wire \w_hssi_gen3_tx_pcs_data_out[1] ;
wire \w_hssi_gen3_tx_pcs_data_out[2] ;
wire \w_hssi_gen3_tx_pcs_data_out[3] ;
wire \w_hssi_gen3_tx_pcs_data_out[4] ;
wire \w_hssi_gen3_tx_pcs_data_out[5] ;
wire \w_hssi_gen3_tx_pcs_data_out[6] ;
wire \w_hssi_gen3_tx_pcs_data_out[7] ;
wire \w_hssi_gen3_tx_pcs_data_out[8] ;
wire \w_hssi_gen3_tx_pcs_data_out[9] ;
wire \w_hssi_gen3_tx_pcs_data_out[10] ;
wire \w_hssi_gen3_tx_pcs_data_out[11] ;
wire \w_hssi_gen3_tx_pcs_data_out[12] ;
wire \w_hssi_gen3_tx_pcs_data_out[13] ;
wire \w_hssi_gen3_tx_pcs_data_out[14] ;
wire \w_hssi_gen3_tx_pcs_data_out[15] ;
wire \w_hssi_gen3_tx_pcs_data_out[16] ;
wire \w_hssi_gen3_tx_pcs_data_out[17] ;
wire \w_hssi_gen3_tx_pcs_data_out[18] ;
wire \w_hssi_gen3_tx_pcs_data_out[19] ;
wire \w_hssi_gen3_tx_pcs_data_out[20] ;
wire \w_hssi_gen3_tx_pcs_data_out[21] ;
wire \w_hssi_gen3_tx_pcs_data_out[22] ;
wire \w_hssi_gen3_tx_pcs_data_out[23] ;
wire \w_hssi_gen3_tx_pcs_data_out[24] ;
wire \w_hssi_gen3_tx_pcs_data_out[25] ;
wire \w_hssi_gen3_tx_pcs_data_out[26] ;
wire \w_hssi_gen3_tx_pcs_data_out[27] ;
wire \w_hssi_gen3_tx_pcs_data_out[28] ;
wire \w_hssi_gen3_tx_pcs_data_out[29] ;
wire \w_hssi_gen3_tx_pcs_data_out[30] ;
wire \w_hssi_gen3_tx_pcs_data_out[31] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[0] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[1] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[2] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[3] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[4] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[5] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[6] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[7] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[8] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[9] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[10] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[11] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[12] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[13] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[14] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[15] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[16] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[17] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[18] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[19] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[20] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[21] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[22] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[23] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[24] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[25] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[26] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[27] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[28] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[29] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[30] ;
wire \w_hssi_gen3_tx_pcs_par_lpbk_out[31] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[0] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[1] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[2] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[3] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[4] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[5] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[6] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[7] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[8] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[9] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[10] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[11] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[12] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[13] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[14] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[15] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[16] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[17] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[18] ;
wire \w_hssi_gen3_tx_pcs_tx_test_out[19] ;
wire w_hssi_krfec_tx_pcs_tx_alignment;
wire w_hssi_krfec_tx_pcs_tx_frame;
wire \w_hssi_krfec_tx_pcs_tx_data_out[0] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[1] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[2] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[3] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[4] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[5] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[6] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[7] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[8] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[9] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[10] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[11] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[12] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[13] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[14] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[15] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[16] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[17] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[18] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[19] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[20] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[21] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[22] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[23] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[24] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[25] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[26] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[27] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[28] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[29] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[30] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[31] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[32] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[33] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[34] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[35] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[36] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[37] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[38] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[39] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[40] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[41] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[42] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[43] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[44] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[45] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[46] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[47] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[48] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[49] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[50] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[51] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[52] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[53] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[54] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[55] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[56] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[57] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[58] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[59] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[60] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[61] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[62] ;
wire \w_hssi_krfec_tx_pcs_tx_data_out[63] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[0] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[1] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[2] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[3] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[4] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[5] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[6] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[7] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[8] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[9] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[10] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[11] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[12] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[13] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[14] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[15] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[16] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[17] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[18] ;
wire \w_hssi_krfec_tx_pcs_tx_test_data[19] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[0] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[1] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[2] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[3] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[4] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[5] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[6] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[7] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[8] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[9] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[10] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[11] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[12] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[13] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[14] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[15] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[16] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[17] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[18] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[19] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[20] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[21] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[22] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[23] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[24] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[25] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[26] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[27] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[28] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[29] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[30] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[31] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[32] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[33] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[34] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[35] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[36] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[37] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[38] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[39] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[40] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[41] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[42] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[43] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[44] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[45] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[46] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[47] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[48] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[49] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[50] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[51] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[52] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[53] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[54] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[55] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[56] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[57] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[58] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[59] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[60] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[61] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[62] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[63] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[64] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[65] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[66] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[67] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[68] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[69] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[70] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[71] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[72] ;
wire \w_hssi_fifo_rx_pcs_data_out2_10g[73] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30] ;
wire \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[0] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[1] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[2] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[3] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[4] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[5] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[6] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[7] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[8] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[9] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[10] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[11] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[12] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[13] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[14] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[15] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[16] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[17] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[18] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[19] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[20] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[21] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[22] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[23] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[24] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[25] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[26] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[27] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[28] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[29] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[30] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[31] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[32] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[33] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[34] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[35] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[36] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[37] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[38] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[39] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[40] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[41] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[42] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[43] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[44] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[45] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[46] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[47] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[48] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[49] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[50] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[51] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[52] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[53] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[54] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[55] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[56] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[57] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[58] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[59] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[60] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[61] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[62] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[63] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[64] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[65] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[66] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[67] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[68] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[69] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[70] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[71] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[72] ;
wire \w_hssi_fifo_rx_pcs_data_out_10g[73] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78] ;
wire \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[0] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[1] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[2] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[3] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[4] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[5] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[6] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[7] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[8] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[9] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[10] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[11] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[12] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[13] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[14] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[15] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[16] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[17] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[18] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[19] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[20] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[21] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[22] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[23] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[24] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[25] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[26] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[27] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[28] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[29] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[30] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[31] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[32] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[33] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[34] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[35] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[36] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[37] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[38] ;
wire \w_hssi_fifo_rx_pcs_data_out_gen3[39] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[0] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[1] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[2] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[3] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[4] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[5] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[6] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[7] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[8] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[9] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[10] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[11] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[12] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[13] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[14] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[15] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[16] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[17] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[18] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[19] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[20] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[21] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[22] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[23] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[24] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[25] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[26] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[27] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[28] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[29] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[30] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[31] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[32] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[33] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[34] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[35] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[36] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[37] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[38] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[39] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[40] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[41] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[42] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[43] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[44] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[45] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[46] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[47] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[48] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[49] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[50] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[51] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[52] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[53] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[54] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[55] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[56] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[57] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[58] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[59] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[60] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[61] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[62] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[63] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[64] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[65] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[66] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[67] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[68] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[69] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[70] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[71] ;
wire \w_hssi_fifo_tx_pcs_data_out_10g[72] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62] ;
wire \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63] ;
wire w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected;
wire w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid;
wire w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done;
wire w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel;
wire w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref;
wire w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6] ;
wire \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7] ;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out;
wire w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out;
wire \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0] ;
wire \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1] ;
wire \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2] ;
wire \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3] ;
wire \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62] ;
wire \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18] ;
wire \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18] ;
wire \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19] ;

wire [7:0] \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus ;
wire [4:0] \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus ;
wire [19:0] \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus ;
wire [127:0] \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus ;
wire [127:0] \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus ;
wire [7:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus ;
wire [2:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_8G_EIDLEINFERSEL_bus ;
wire [17:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus ;
wire [2:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_RXPRESET_bus ;
wire [5:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus ;
wire [1:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PCIE_SWITCH_bus ;
wire [4:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus ;
wire [1:0] \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_RATE_bus ;
wire [7:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus ;
wire [6:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus ;
wire [17:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus ;
wire [8:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus ;
wire [127:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus ;
wire [1:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DIAG_STATUS_bus ;
wire [1:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_POWERDOWN_bus ;
wire [3:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus ;
wire [4:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus ;
wire [3:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus ;
wire [1:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_SYNC_HDR_bus ;
wire [43:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus ;
wire [43:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus ;
wire [2:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXMARGIN_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus ;
wire [19:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus ;
wire [127:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus ;
wire [7:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus ;
wire [1:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DIAG_STATUS_bus ;
wire [4:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus ;
wire [31:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus ;
wire [31:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus ;
wire [73:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus ;
wire [31:0] \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus ;
wire [4:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus ;
wire [19:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus ;
wire [63:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus ;
wire [3:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus ;
wire [7:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus ;
wire [63:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus ;
wire [3:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus ;
wire [2:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RXSTATUS_bus ;
wire [19:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus ;
wire [2:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_EIOS_DET_CDR_CTRL_bus ;
wire [19:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus ;
wire [19:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus ;
wire [7:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus ;
wire [3:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus ;
wire [1:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_SYNC_HDR_bus ;
wire [79:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus ;
wire [31:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus ;
wire [7:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus ;
wire [19:0] \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus ;
wire [7:0] \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus ;
wire [2:0] \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_RXSTATUS_bus ;
wire [17:0] \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus ;
wire [7:0] \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus ;
wire [9:0] \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus ;
wire [63:0] \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus ;
wire [1:0] \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_STATUS_bus ;
wire [7:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus ;
wire [63:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus ;
wire [19:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus ;
wire [31:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus ;
wire [63:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus ;
wire [5:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus ;
wire [19:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus ;
wire [19:0] \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus ;
wire [7:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus ;
wire [19:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus ;
wire [2:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_NON_GRAY_EIDLEINFERSEL_bus ;
wire [2:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PHFIFO_TXMARGIN_bus ;
wire [7:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus ;
wire [3:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_BLK_START_OUT_bus ;
wire [19:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus ;
wire [31:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus ;
wire [3:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_VALID_OUT_bus ;
wire [3:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus ;
wire [1:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DIV_SYNC_bus ;
wire [1:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_SYNC_HDR_OUT_bus ;
wire [19:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus ;
wire [63:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus ;
wire [7:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus ;
wire [1:0] \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PIPE_POWER_DOWN_OUT_bus ;
wire [63:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus ;
wire [7:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus ;
wire [8:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus ;
wire [63:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus ;
wire [3:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus ;
wire [15:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus ;
wire [72:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus ;
wire [72:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus ;
wire [15:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus ;
wire [63:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus ;
wire [19:0] \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus ;
wire [31:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus ;
wire [33:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus ;
wire [15:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus ;
wire [39:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus ;
wire [15:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus ;
wire [19:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus ;
wire [1:0] \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_SYNC_HDR_bus ;
wire [19:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus ;
wire [2:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXSTATUS_bus ;
wire [3:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus ;
wire [1:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_SYNC_HDR_bus ;
wire [17:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus ;
wire [2:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_RXPRESET_bus ;
wire [63:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus ;
wire [3:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus ;
wire [1:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TX_SYNC_HDR_INT_bus ;
wire [31:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus ;
wire [3:0] \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus ;
wire [31:0] \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus ;
wire [35:0] \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus ;
wire [31:0] \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus ;
wire [19:0] \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus ;
wire [19:0] \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus ;
wire [73:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus ;
wire [31:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus ;
wire [73:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus ;
wire [31:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus ;
wire [79:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus ;
wire [39:0] \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus ;
wire [7:0] \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus ;
wire [72:0] \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus ;
wire [63:0] \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus ;
wire [7:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus ;
wire [8:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus ;
wire [8:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus ;
wire [1:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PCIE_SW_DONE_bus ;
wire [4:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus ;
wire [19:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus ;
wire [7:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus ;
wire [17:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus ;
wire [1:0] \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_PCIE_SWITCH_bus ;
wire [7:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus ;
wire [15:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus ;
wire [4:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus ;
wire [63:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus ;
wire [19:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus ;
wire [19:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus ;
wire [19:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus ;
wire [19:0] \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus ;

assign out_avmmreaddata_hssi_rx_pld_pcs_interface[0] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[1] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[2] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[3] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[4] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[5] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[6] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_rx_pld_pcs_interface[7] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus [7];

assign out_pld_8g_wa_boundary[0] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus [0];
assign out_pld_8g_wa_boundary[1] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus [1];
assign out_pld_8g_wa_boundary[2] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus [2];
assign out_pld_8g_wa_boundary[3] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus [3];
assign out_pld_8g_wa_boundary[4] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus [4];

assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [0];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [1];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [2];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [3];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [4];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [5];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [6];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [7];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [8];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [9];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [10];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [11];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [12];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [13];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [14];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [15];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [16];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [17];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [18];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus [19];

assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [0];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [1];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [2];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [3];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [4];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [5];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [6];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [7];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [8];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [9];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [10];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [11];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [12];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [13];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [14];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [15];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [16];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [17];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [18];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [19];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [20];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [21];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [22];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [23];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [24];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [25];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [26];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [27];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [28];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [29];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [30];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [31];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [32];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [33];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [34];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [35];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [36];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [37];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [38];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [39];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [40];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [41];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [42];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [43];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [44];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [45];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [46];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [47];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [48];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [49];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [50];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [51];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [52];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [53];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [54];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [55];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [56];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [57];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [58];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [59];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [60];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [61];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [62];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [63];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [64];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [65];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [66];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [67];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [68];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [69];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [70];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [71];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [72];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [73];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [74];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [75];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [76];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [77];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [78];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [79];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [80];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [81];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [82];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [83];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [84];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [85];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [86];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [87];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [88];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [89];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [90];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [91];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [92];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [93];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [94];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [95];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [96];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [97];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [98];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [99];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [100];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [101];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [102];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [103];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [104];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [105];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [106];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [107];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [108];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [109];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [110];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [111];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [112];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [113];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [114];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [115];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [116];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [117];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [118];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [119];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [120];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [121];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [122];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [123];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [124];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [125];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [126];
assign \w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127]  = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus [127];

assign out_pld_rx_data[0] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [0];
assign out_pld_rx_data[1] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [1];
assign out_pld_rx_data[2] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [2];
assign out_pld_rx_data[3] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [3];
assign out_pld_rx_data[4] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [4];
assign out_pld_rx_data[5] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [5];
assign out_pld_rx_data[6] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [6];
assign out_pld_rx_data[7] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [7];
assign out_pld_rx_data[8] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [8];
assign out_pld_rx_data[9] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [9];
assign out_pld_rx_data[10] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [10];
assign out_pld_rx_data[11] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [11];
assign out_pld_rx_data[12] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [12];
assign out_pld_rx_data[13] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [13];
assign out_pld_rx_data[14] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [14];
assign out_pld_rx_data[15] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [15];
assign out_pld_rx_data[16] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [16];
assign out_pld_rx_data[17] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [17];
assign out_pld_rx_data[18] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [18];
assign out_pld_rx_data[19] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [19];
assign out_pld_rx_data[20] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [20];
assign out_pld_rx_data[21] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [21];
assign out_pld_rx_data[22] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [22];
assign out_pld_rx_data[23] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [23];
assign out_pld_rx_data[24] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [24];
assign out_pld_rx_data[25] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [25];
assign out_pld_rx_data[26] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [26];
assign out_pld_rx_data[27] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [27];
assign out_pld_rx_data[28] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [28];
assign out_pld_rx_data[29] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [29];
assign out_pld_rx_data[30] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [30];
assign out_pld_rx_data[31] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [31];
assign out_pld_rx_data[32] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [32];
assign out_pld_rx_data[33] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [33];
assign out_pld_rx_data[34] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [34];
assign out_pld_rx_data[35] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [35];
assign out_pld_rx_data[36] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [36];
assign out_pld_rx_data[37] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [37];
assign out_pld_rx_data[38] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [38];
assign out_pld_rx_data[39] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [39];
assign out_pld_rx_data[40] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [40];
assign out_pld_rx_data[41] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [41];
assign out_pld_rx_data[42] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [42];
assign out_pld_rx_data[43] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [43];
assign out_pld_rx_data[44] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [44];
assign out_pld_rx_data[45] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [45];
assign out_pld_rx_data[46] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [46];
assign out_pld_rx_data[47] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [47];
assign out_pld_rx_data[48] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [48];
assign out_pld_rx_data[49] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [49];
assign out_pld_rx_data[50] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [50];
assign out_pld_rx_data[51] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [51];
assign out_pld_rx_data[52] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [52];
assign out_pld_rx_data[53] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [53];
assign out_pld_rx_data[54] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [54];
assign out_pld_rx_data[55] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [55];
assign out_pld_rx_data[56] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [56];
assign out_pld_rx_data[57] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [57];
assign out_pld_rx_data[58] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [58];
assign out_pld_rx_data[59] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [59];
assign out_pld_rx_data[60] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [60];
assign out_pld_rx_data[61] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [61];
assign out_pld_rx_data[62] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [62];
assign out_pld_rx_data[63] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [63];
assign out_pld_rx_data[64] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [64];
assign out_pld_rx_data[65] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [65];
assign out_pld_rx_data[66] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [66];
assign out_pld_rx_data[67] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [67];
assign out_pld_rx_data[68] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [68];
assign out_pld_rx_data[69] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [69];
assign out_pld_rx_data[70] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [70];
assign out_pld_rx_data[71] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [71];
assign out_pld_rx_data[72] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [72];
assign out_pld_rx_data[73] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [73];
assign out_pld_rx_data[74] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [74];
assign out_pld_rx_data[75] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [75];
assign out_pld_rx_data[76] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [76];
assign out_pld_rx_data[77] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [77];
assign out_pld_rx_data[78] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [78];
assign out_pld_rx_data[79] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [79];
assign out_pld_rx_data[80] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [80];
assign out_pld_rx_data[81] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [81];
assign out_pld_rx_data[82] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [82];
assign out_pld_rx_data[83] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [83];
assign out_pld_rx_data[84] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [84];
assign out_pld_rx_data[85] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [85];
assign out_pld_rx_data[86] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [86];
assign out_pld_rx_data[87] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [87];
assign out_pld_rx_data[88] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [88];
assign out_pld_rx_data[89] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [89];
assign out_pld_rx_data[90] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [90];
assign out_pld_rx_data[91] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [91];
assign out_pld_rx_data[92] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [92];
assign out_pld_rx_data[93] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [93];
assign out_pld_rx_data[94] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [94];
assign out_pld_rx_data[95] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [95];
assign out_pld_rx_data[96] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [96];
assign out_pld_rx_data[97] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [97];
assign out_pld_rx_data[98] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [98];
assign out_pld_rx_data[99] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [99];
assign out_pld_rx_data[100] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [100];
assign out_pld_rx_data[101] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [101];
assign out_pld_rx_data[102] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [102];
assign out_pld_rx_data[103] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [103];
assign out_pld_rx_data[104] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [104];
assign out_pld_rx_data[105] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [105];
assign out_pld_rx_data[106] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [106];
assign out_pld_rx_data[107] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [107];
assign out_pld_rx_data[108] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [108];
assign out_pld_rx_data[109] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [109];
assign out_pld_rx_data[110] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [110];
assign out_pld_rx_data[111] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [111];
assign out_pld_rx_data[112] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [112];
assign out_pld_rx_data[113] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [113];
assign out_pld_rx_data[114] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [114];
assign out_pld_rx_data[115] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [115];
assign out_pld_rx_data[116] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [116];
assign out_pld_rx_data[117] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [117];
assign out_pld_rx_data[118] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [118];
assign out_pld_rx_data[119] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [119];
assign out_pld_rx_data[120] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [120];
assign out_pld_rx_data[121] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [121];
assign out_pld_rx_data[122] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [122];
assign out_pld_rx_data[123] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [123];
assign out_pld_rx_data[124] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [124];
assign out_pld_rx_data[125] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [125];
assign out_pld_rx_data[126] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [126];
assign out_pld_rx_data[127] = \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus [127];

assign out_avmmreaddata_hssi_common_pld_pcs_interface[0] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[1] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[2] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[3] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[4] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[5] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[6] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_common_pld_pcs_interface[7] = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus [7];

assign \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_8G_EIDLEINFERSEL_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_8G_EIDLEINFERSEL_bus [1];
assign \w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_8G_EIDLEINFERSEL_bus [2];

assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [1];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [2];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [3];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [4];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [5];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [6];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [7];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [8];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [9];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [10];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [11];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [12];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [13];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [14];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [15];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [16];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus [17];

assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_RXPRESET_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_RXPRESET_bus [1];
assign \w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_RXPRESET_bus [2];

assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [1];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [2];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [3];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [4];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus [5];

assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PCIE_SWITCH_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PCIE_SWITCH_bus [1];

assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus [1];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus [2];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus [3];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus [4];

assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_RATE_bus [0];
assign \w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1]  = \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_RATE_bus [1];

assign out_avmmreaddata_hssi_tx_pld_pcs_interface[0] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[1] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[2] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[3] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[4] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[5] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[6] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_tx_pld_pcs_interface[7] = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus [7];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus [6];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus [17];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus [8];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [43];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [44];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [45];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [46];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [47];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [48];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [49];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [50];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [51];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [52];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [53];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [54];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [55];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [56];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [57];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [58];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [59];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [60];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [61];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [62];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [63];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [64];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [65];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [66];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [67];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [68];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [69];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [70];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [71];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [72];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [73];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [74];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [75];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [76];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [77];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [78];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [79];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [80];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [81];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [82];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [83];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [84];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [85];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [86];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [87];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [88];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [89];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [90];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [91];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [92];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [93];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [94];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [95];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [96];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [97];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [98];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [99];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [100];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [101];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [102];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [103];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [104];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [105];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [106];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [107];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [108];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [109];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [110];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [111];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [112];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [113];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [114];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [115];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [116];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [117];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [118];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [119];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [120];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [121];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [122];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [123];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [124];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [125];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [126];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus [127];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [43];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [44];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [45];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [46];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [47];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [48];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [49];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [50];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [51];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [52];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [53];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [54];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [55];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [56];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [57];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [58];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [59];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [60];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [61];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [62];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus [63];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DIAG_STATUS_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DIAG_STATUS_bus [1];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_POWERDOWN_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_POWERDOWN_bus [1];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus [3];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus [4];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus [3];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_SYNC_HDR_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_SYNC_HDR_bus [1];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus [43];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus [43];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXMARGIN_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXMARGIN_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXMARGIN_bus [2];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [43];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [44];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [45];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [46];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [47];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [48];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [49];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [50];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [51];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [52];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [53];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [54];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [55];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [56];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [57];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [58];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [59];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [60];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [61];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [62];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus [63];

assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [0];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [1];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [2];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [3];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [4];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [5];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [6];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [7];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [8];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [9];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [10];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [11];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [12];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [13];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [14];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [15];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [16];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [17];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [18];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [19];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [20];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [21];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [22];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [23];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [24];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [25];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [26];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [27];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [28];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [29];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [30];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [31];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [32];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [33];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [34];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [35];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [36];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [37];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [38];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [39];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [40];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [41];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [42];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [43];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [44];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [45];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [46];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [47];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [48];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [49];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [50];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [51];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [52];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [53];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [54];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [55];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [56];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [57];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [58];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [59];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [60];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [61];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [62];
assign \w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63]  = \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus [63];

assign \w_hssi_10g_rx_pcs_rx_control[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [0];
assign \w_hssi_10g_rx_pcs_rx_control[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [1];
assign \w_hssi_10g_rx_pcs_rx_control[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [2];
assign \w_hssi_10g_rx_pcs_rx_control[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [3];
assign \w_hssi_10g_rx_pcs_rx_control[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [4];
assign \w_hssi_10g_rx_pcs_rx_control[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [5];
assign \w_hssi_10g_rx_pcs_rx_control[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [6];
assign \w_hssi_10g_rx_pcs_rx_control[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [7];
assign \w_hssi_10g_rx_pcs_rx_control[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [8];
assign \w_hssi_10g_rx_pcs_rx_control[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [9];
assign \w_hssi_10g_rx_pcs_rx_control[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [10];
assign \w_hssi_10g_rx_pcs_rx_control[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [11];
assign \w_hssi_10g_rx_pcs_rx_control[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [12];
assign \w_hssi_10g_rx_pcs_rx_control[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [13];
assign \w_hssi_10g_rx_pcs_rx_control[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [14];
assign \w_hssi_10g_rx_pcs_rx_control[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [15];
assign \w_hssi_10g_rx_pcs_rx_control[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [16];
assign \w_hssi_10g_rx_pcs_rx_control[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [17];
assign \w_hssi_10g_rx_pcs_rx_control[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [18];
assign \w_hssi_10g_rx_pcs_rx_control[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus [19];

assign \w_hssi_10g_rx_pcs_rx_data[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [0];
assign \w_hssi_10g_rx_pcs_rx_data[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [1];
assign \w_hssi_10g_rx_pcs_rx_data[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [2];
assign \w_hssi_10g_rx_pcs_rx_data[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [3];
assign \w_hssi_10g_rx_pcs_rx_data[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [4];
assign \w_hssi_10g_rx_pcs_rx_data[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [5];
assign \w_hssi_10g_rx_pcs_rx_data[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [6];
assign \w_hssi_10g_rx_pcs_rx_data[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [7];
assign \w_hssi_10g_rx_pcs_rx_data[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [8];
assign \w_hssi_10g_rx_pcs_rx_data[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [9];
assign \w_hssi_10g_rx_pcs_rx_data[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [10];
assign \w_hssi_10g_rx_pcs_rx_data[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [11];
assign \w_hssi_10g_rx_pcs_rx_data[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [12];
assign \w_hssi_10g_rx_pcs_rx_data[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [13];
assign \w_hssi_10g_rx_pcs_rx_data[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [14];
assign \w_hssi_10g_rx_pcs_rx_data[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [15];
assign \w_hssi_10g_rx_pcs_rx_data[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [16];
assign \w_hssi_10g_rx_pcs_rx_data[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [17];
assign \w_hssi_10g_rx_pcs_rx_data[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [18];
assign \w_hssi_10g_rx_pcs_rx_data[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [19];
assign \w_hssi_10g_rx_pcs_rx_data[20]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [20];
assign \w_hssi_10g_rx_pcs_rx_data[21]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [21];
assign \w_hssi_10g_rx_pcs_rx_data[22]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [22];
assign \w_hssi_10g_rx_pcs_rx_data[23]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [23];
assign \w_hssi_10g_rx_pcs_rx_data[24]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [24];
assign \w_hssi_10g_rx_pcs_rx_data[25]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [25];
assign \w_hssi_10g_rx_pcs_rx_data[26]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [26];
assign \w_hssi_10g_rx_pcs_rx_data[27]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [27];
assign \w_hssi_10g_rx_pcs_rx_data[28]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [28];
assign \w_hssi_10g_rx_pcs_rx_data[29]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [29];
assign \w_hssi_10g_rx_pcs_rx_data[30]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [30];
assign \w_hssi_10g_rx_pcs_rx_data[31]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [31];
assign \w_hssi_10g_rx_pcs_rx_data[32]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [32];
assign \w_hssi_10g_rx_pcs_rx_data[33]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [33];
assign \w_hssi_10g_rx_pcs_rx_data[34]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [34];
assign \w_hssi_10g_rx_pcs_rx_data[35]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [35];
assign \w_hssi_10g_rx_pcs_rx_data[36]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [36];
assign \w_hssi_10g_rx_pcs_rx_data[37]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [37];
assign \w_hssi_10g_rx_pcs_rx_data[38]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [38];
assign \w_hssi_10g_rx_pcs_rx_data[39]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [39];
assign \w_hssi_10g_rx_pcs_rx_data[40]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [40];
assign \w_hssi_10g_rx_pcs_rx_data[41]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [41];
assign \w_hssi_10g_rx_pcs_rx_data[42]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [42];
assign \w_hssi_10g_rx_pcs_rx_data[43]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [43];
assign \w_hssi_10g_rx_pcs_rx_data[44]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [44];
assign \w_hssi_10g_rx_pcs_rx_data[45]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [45];
assign \w_hssi_10g_rx_pcs_rx_data[46]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [46];
assign \w_hssi_10g_rx_pcs_rx_data[47]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [47];
assign \w_hssi_10g_rx_pcs_rx_data[48]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [48];
assign \w_hssi_10g_rx_pcs_rx_data[49]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [49];
assign \w_hssi_10g_rx_pcs_rx_data[50]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [50];
assign \w_hssi_10g_rx_pcs_rx_data[51]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [51];
assign \w_hssi_10g_rx_pcs_rx_data[52]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [52];
assign \w_hssi_10g_rx_pcs_rx_data[53]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [53];
assign \w_hssi_10g_rx_pcs_rx_data[54]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [54];
assign \w_hssi_10g_rx_pcs_rx_data[55]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [55];
assign \w_hssi_10g_rx_pcs_rx_data[56]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [56];
assign \w_hssi_10g_rx_pcs_rx_data[57]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [57];
assign \w_hssi_10g_rx_pcs_rx_data[58]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [58];
assign \w_hssi_10g_rx_pcs_rx_data[59]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [59];
assign \w_hssi_10g_rx_pcs_rx_data[60]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [60];
assign \w_hssi_10g_rx_pcs_rx_data[61]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [61];
assign \w_hssi_10g_rx_pcs_rx_data[62]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [62];
assign \w_hssi_10g_rx_pcs_rx_data[63]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [63];
assign \w_hssi_10g_rx_pcs_rx_data[64]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [64];
assign \w_hssi_10g_rx_pcs_rx_data[65]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [65];
assign \w_hssi_10g_rx_pcs_rx_data[66]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [66];
assign \w_hssi_10g_rx_pcs_rx_data[67]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [67];
assign \w_hssi_10g_rx_pcs_rx_data[68]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [68];
assign \w_hssi_10g_rx_pcs_rx_data[69]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [69];
assign \w_hssi_10g_rx_pcs_rx_data[70]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [70];
assign \w_hssi_10g_rx_pcs_rx_data[71]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [71];
assign \w_hssi_10g_rx_pcs_rx_data[72]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [72];
assign \w_hssi_10g_rx_pcs_rx_data[73]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [73];
assign \w_hssi_10g_rx_pcs_rx_data[74]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [74];
assign \w_hssi_10g_rx_pcs_rx_data[75]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [75];
assign \w_hssi_10g_rx_pcs_rx_data[76]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [76];
assign \w_hssi_10g_rx_pcs_rx_data[77]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [77];
assign \w_hssi_10g_rx_pcs_rx_data[78]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [78];
assign \w_hssi_10g_rx_pcs_rx_data[79]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [79];
assign \w_hssi_10g_rx_pcs_rx_data[80]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [80];
assign \w_hssi_10g_rx_pcs_rx_data[81]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [81];
assign \w_hssi_10g_rx_pcs_rx_data[82]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [82];
assign \w_hssi_10g_rx_pcs_rx_data[83]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [83];
assign \w_hssi_10g_rx_pcs_rx_data[84]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [84];
assign \w_hssi_10g_rx_pcs_rx_data[85]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [85];
assign \w_hssi_10g_rx_pcs_rx_data[86]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [86];
assign \w_hssi_10g_rx_pcs_rx_data[87]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [87];
assign \w_hssi_10g_rx_pcs_rx_data[88]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [88];
assign \w_hssi_10g_rx_pcs_rx_data[89]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [89];
assign \w_hssi_10g_rx_pcs_rx_data[90]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [90];
assign \w_hssi_10g_rx_pcs_rx_data[91]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [91];
assign \w_hssi_10g_rx_pcs_rx_data[92]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [92];
assign \w_hssi_10g_rx_pcs_rx_data[93]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [93];
assign \w_hssi_10g_rx_pcs_rx_data[94]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [94];
assign \w_hssi_10g_rx_pcs_rx_data[95]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [95];
assign \w_hssi_10g_rx_pcs_rx_data[96]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [96];
assign \w_hssi_10g_rx_pcs_rx_data[97]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [97];
assign \w_hssi_10g_rx_pcs_rx_data[98]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [98];
assign \w_hssi_10g_rx_pcs_rx_data[99]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [99];
assign \w_hssi_10g_rx_pcs_rx_data[100]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [100];
assign \w_hssi_10g_rx_pcs_rx_data[101]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [101];
assign \w_hssi_10g_rx_pcs_rx_data[102]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [102];
assign \w_hssi_10g_rx_pcs_rx_data[103]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [103];
assign \w_hssi_10g_rx_pcs_rx_data[104]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [104];
assign \w_hssi_10g_rx_pcs_rx_data[105]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [105];
assign \w_hssi_10g_rx_pcs_rx_data[106]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [106];
assign \w_hssi_10g_rx_pcs_rx_data[107]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [107];
assign \w_hssi_10g_rx_pcs_rx_data[108]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [108];
assign \w_hssi_10g_rx_pcs_rx_data[109]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [109];
assign \w_hssi_10g_rx_pcs_rx_data[110]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [110];
assign \w_hssi_10g_rx_pcs_rx_data[111]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [111];
assign \w_hssi_10g_rx_pcs_rx_data[112]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [112];
assign \w_hssi_10g_rx_pcs_rx_data[113]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [113];
assign \w_hssi_10g_rx_pcs_rx_data[114]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [114];
assign \w_hssi_10g_rx_pcs_rx_data[115]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [115];
assign \w_hssi_10g_rx_pcs_rx_data[116]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [116];
assign \w_hssi_10g_rx_pcs_rx_data[117]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [117];
assign \w_hssi_10g_rx_pcs_rx_data[118]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [118];
assign \w_hssi_10g_rx_pcs_rx_data[119]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [119];
assign \w_hssi_10g_rx_pcs_rx_data[120]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [120];
assign \w_hssi_10g_rx_pcs_rx_data[121]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [121];
assign \w_hssi_10g_rx_pcs_rx_data[122]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [122];
assign \w_hssi_10g_rx_pcs_rx_data[123]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [123];
assign \w_hssi_10g_rx_pcs_rx_data[124]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [124];
assign \w_hssi_10g_rx_pcs_rx_data[125]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [125];
assign \w_hssi_10g_rx_pcs_rx_data[126]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [126];
assign \w_hssi_10g_rx_pcs_rx_data[127]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus [127];

assign out_avmmreaddata_hssi_10g_rx_pcs[0] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_10g_rx_pcs[1] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_10g_rx_pcs[2] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_10g_rx_pcs[3] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_10g_rx_pcs[4] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_10g_rx_pcs[5] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_10g_rx_pcs[6] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_10g_rx_pcs[7] = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_10g_rx_pcs_rx_diag_status[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DIAG_STATUS_bus [0];
assign \w_hssi_10g_rx_pcs_rx_diag_status[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DIAG_STATUS_bus [1];

assign \w_hssi_10g_rx_pcs_rx_fifo_num[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus [0];
assign \w_hssi_10g_rx_pcs_rx_fifo_num[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus [1];
assign \w_hssi_10g_rx_pcs_rx_fifo_num[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus [2];
assign \w_hssi_10g_rx_pcs_rx_fifo_num[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus [3];
assign \w_hssi_10g_rx_pcs_rx_fifo_num[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus [4];

assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [0];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [1];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [2];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [3];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [4];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [5];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [6];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [7];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [8];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [9];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [10];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [11];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [12];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [13];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [14];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [15];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [16];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [17];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [18];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [19];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [20];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [21];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [22];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [23];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [24];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [25];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [26];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [27];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [28];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [29];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [30];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus [31];

assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [0];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [1];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [2];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [3];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [4];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [5];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [6];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [7];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [8];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [9];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [10];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [11];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [12];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [13];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [14];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [15];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [16];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [17];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [18];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [19];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [20];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [21];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [22];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [23];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [24];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [25];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [26];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [27];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [28];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [29];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [30];
assign \w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus [31];

assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [0];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [1];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [2];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [3];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [4];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [5];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [6];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [7];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [8];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [9];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [10];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [11];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [12];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [13];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [14];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [15];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [16];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [17];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [18];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [19];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[20]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [20];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[21]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [21];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[22]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [22];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[23]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [23];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[24]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [24];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[25]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [25];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[26]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [26];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[27]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [27];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[28]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [28];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[29]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [29];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[30]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [30];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[31]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [31];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[32]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [32];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[33]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [33];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[34]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [34];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[35]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [35];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[36]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [36];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[37]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [37];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[38]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [38];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[39]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [39];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[40]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [40];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[41]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [41];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[42]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [42];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[43]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [43];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[44]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [44];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[45]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [45];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[46]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [46];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[47]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [47];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[48]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [48];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[49]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [49];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[50]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [50];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[51]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [51];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[52]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [52];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[53]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [53];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[54]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [54];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[55]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [55];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[56]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [56];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[57]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [57];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[58]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [58];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[59]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [59];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[60]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [60];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[61]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [61];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[62]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [62];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[63]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [63];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[64]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [64];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[65]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [65];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[66]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [66];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[67]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [67];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[68]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [68];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[69]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [69];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[70]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [70];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[71]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [71];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[72]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [72];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_data[73]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus [73];

assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [0];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [1];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [2];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [3];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [4];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [5];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [6];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [7];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [8];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [9];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [10];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [11];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [12];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [13];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [14];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [15];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [16];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [17];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [18];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [19];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [20];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [21];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [22];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [23];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [24];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [25];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [26];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [27];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [28];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [29];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [30];
assign \w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31]  = \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus [31];

assign \w_hssi_8g_rx_pcs_word_align_boundary[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus [0];
assign \w_hssi_8g_rx_pcs_word_align_boundary[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus [1];
assign \w_hssi_8g_rx_pcs_word_align_boundary[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus [2];
assign \w_hssi_8g_rx_pcs_word_align_boundary[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus [3];
assign \w_hssi_8g_rx_pcs_word_align_boundary[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus [4];

assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [0];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [1];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [2];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [3];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [4];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [5];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [6];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [7];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [8];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [9];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [10];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [11];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [12];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [13];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [14];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [15];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [16];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [17];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [18];
assign \w_hssi_8g_rx_pcs_parallel_rev_loopback[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus [19];

assign \w_hssi_8g_rx_pcs_pipe_data[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [0];
assign \w_hssi_8g_rx_pcs_pipe_data[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [1];
assign \w_hssi_8g_rx_pcs_pipe_data[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [2];
assign \w_hssi_8g_rx_pcs_pipe_data[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [3];
assign \w_hssi_8g_rx_pcs_pipe_data[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [4];
assign \w_hssi_8g_rx_pcs_pipe_data[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [5];
assign \w_hssi_8g_rx_pcs_pipe_data[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [6];
assign \w_hssi_8g_rx_pcs_pipe_data[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [7];
assign \w_hssi_8g_rx_pcs_pipe_data[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [8];
assign \w_hssi_8g_rx_pcs_pipe_data[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [9];
assign \w_hssi_8g_rx_pcs_pipe_data[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [10];
assign \w_hssi_8g_rx_pcs_pipe_data[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [11];
assign \w_hssi_8g_rx_pcs_pipe_data[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [12];
assign \w_hssi_8g_rx_pcs_pipe_data[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [13];
assign \w_hssi_8g_rx_pcs_pipe_data[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [14];
assign \w_hssi_8g_rx_pcs_pipe_data[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [15];
assign \w_hssi_8g_rx_pcs_pipe_data[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [16];
assign \w_hssi_8g_rx_pcs_pipe_data[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [17];
assign \w_hssi_8g_rx_pcs_pipe_data[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [18];
assign \w_hssi_8g_rx_pcs_pipe_data[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [19];
assign \w_hssi_8g_rx_pcs_pipe_data[20]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [20];
assign \w_hssi_8g_rx_pcs_pipe_data[21]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [21];
assign \w_hssi_8g_rx_pcs_pipe_data[22]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [22];
assign \w_hssi_8g_rx_pcs_pipe_data[23]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [23];
assign \w_hssi_8g_rx_pcs_pipe_data[24]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [24];
assign \w_hssi_8g_rx_pcs_pipe_data[25]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [25];
assign \w_hssi_8g_rx_pcs_pipe_data[26]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [26];
assign \w_hssi_8g_rx_pcs_pipe_data[27]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [27];
assign \w_hssi_8g_rx_pcs_pipe_data[28]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [28];
assign \w_hssi_8g_rx_pcs_pipe_data[29]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [29];
assign \w_hssi_8g_rx_pcs_pipe_data[30]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [30];
assign \w_hssi_8g_rx_pcs_pipe_data[31]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [31];
assign \w_hssi_8g_rx_pcs_pipe_data[32]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [32];
assign \w_hssi_8g_rx_pcs_pipe_data[33]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [33];
assign \w_hssi_8g_rx_pcs_pipe_data[34]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [34];
assign \w_hssi_8g_rx_pcs_pipe_data[35]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [35];
assign \w_hssi_8g_rx_pcs_pipe_data[36]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [36];
assign \w_hssi_8g_rx_pcs_pipe_data[37]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [37];
assign \w_hssi_8g_rx_pcs_pipe_data[38]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [38];
assign \w_hssi_8g_rx_pcs_pipe_data[39]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [39];
assign \w_hssi_8g_rx_pcs_pipe_data[40]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [40];
assign \w_hssi_8g_rx_pcs_pipe_data[41]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [41];
assign \w_hssi_8g_rx_pcs_pipe_data[42]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [42];
assign \w_hssi_8g_rx_pcs_pipe_data[43]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [43];
assign \w_hssi_8g_rx_pcs_pipe_data[44]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [44];
assign \w_hssi_8g_rx_pcs_pipe_data[45]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [45];
assign \w_hssi_8g_rx_pcs_pipe_data[46]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [46];
assign \w_hssi_8g_rx_pcs_pipe_data[47]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [47];
assign \w_hssi_8g_rx_pcs_pipe_data[48]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [48];
assign \w_hssi_8g_rx_pcs_pipe_data[49]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [49];
assign \w_hssi_8g_rx_pcs_pipe_data[50]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [50];
assign \w_hssi_8g_rx_pcs_pipe_data[51]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [51];
assign \w_hssi_8g_rx_pcs_pipe_data[52]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [52];
assign \w_hssi_8g_rx_pcs_pipe_data[53]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [53];
assign \w_hssi_8g_rx_pcs_pipe_data[54]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [54];
assign \w_hssi_8g_rx_pcs_pipe_data[55]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [55];
assign \w_hssi_8g_rx_pcs_pipe_data[56]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [56];
assign \w_hssi_8g_rx_pcs_pipe_data[57]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [57];
assign \w_hssi_8g_rx_pcs_pipe_data[58]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [58];
assign \w_hssi_8g_rx_pcs_pipe_data[59]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [59];
assign \w_hssi_8g_rx_pcs_pipe_data[60]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [60];
assign \w_hssi_8g_rx_pcs_pipe_data[61]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [61];
assign \w_hssi_8g_rx_pcs_pipe_data[62]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [62];
assign \w_hssi_8g_rx_pcs_pipe_data[63]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus [63];

assign \w_hssi_8g_rx_pcs_rx_data_valid[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus [0];
assign \w_hssi_8g_rx_pcs_rx_data_valid[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus [1];
assign \w_hssi_8g_rx_pcs_rx_data_valid[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus [2];
assign \w_hssi_8g_rx_pcs_rx_data_valid[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus [3];

assign out_avmmreaddata_hssi_8g_rx_pcs[0] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_8g_rx_pcs[1] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_8g_rx_pcs[2] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_8g_rx_pcs[3] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_8g_rx_pcs[4] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_8g_rx_pcs[5] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_8g_rx_pcs[6] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_8g_rx_pcs[7] = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_8g_rx_pcs_dataout[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [0];
assign \w_hssi_8g_rx_pcs_dataout[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [1];
assign \w_hssi_8g_rx_pcs_dataout[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [2];
assign \w_hssi_8g_rx_pcs_dataout[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [3];
assign \w_hssi_8g_rx_pcs_dataout[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [4];
assign \w_hssi_8g_rx_pcs_dataout[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [5];
assign \w_hssi_8g_rx_pcs_dataout[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [6];
assign \w_hssi_8g_rx_pcs_dataout[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [7];
assign \w_hssi_8g_rx_pcs_dataout[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [8];
assign \w_hssi_8g_rx_pcs_dataout[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [9];
assign \w_hssi_8g_rx_pcs_dataout[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [10];
assign \w_hssi_8g_rx_pcs_dataout[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [11];
assign \w_hssi_8g_rx_pcs_dataout[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [12];
assign \w_hssi_8g_rx_pcs_dataout[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [13];
assign \w_hssi_8g_rx_pcs_dataout[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [14];
assign \w_hssi_8g_rx_pcs_dataout[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [15];
assign \w_hssi_8g_rx_pcs_dataout[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [16];
assign \w_hssi_8g_rx_pcs_dataout[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [17];
assign \w_hssi_8g_rx_pcs_dataout[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [18];
assign \w_hssi_8g_rx_pcs_dataout[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [19];
assign \w_hssi_8g_rx_pcs_dataout[20]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [20];
assign \w_hssi_8g_rx_pcs_dataout[21]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [21];
assign \w_hssi_8g_rx_pcs_dataout[22]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [22];
assign \w_hssi_8g_rx_pcs_dataout[23]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [23];
assign \w_hssi_8g_rx_pcs_dataout[24]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [24];
assign \w_hssi_8g_rx_pcs_dataout[25]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [25];
assign \w_hssi_8g_rx_pcs_dataout[26]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [26];
assign \w_hssi_8g_rx_pcs_dataout[27]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [27];
assign \w_hssi_8g_rx_pcs_dataout[28]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [28];
assign \w_hssi_8g_rx_pcs_dataout[29]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [29];
assign \w_hssi_8g_rx_pcs_dataout[30]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [30];
assign \w_hssi_8g_rx_pcs_dataout[31]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [31];
assign \w_hssi_8g_rx_pcs_dataout[32]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [32];
assign \w_hssi_8g_rx_pcs_dataout[33]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [33];
assign \w_hssi_8g_rx_pcs_dataout[34]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [34];
assign \w_hssi_8g_rx_pcs_dataout[35]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [35];
assign \w_hssi_8g_rx_pcs_dataout[36]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [36];
assign \w_hssi_8g_rx_pcs_dataout[37]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [37];
assign \w_hssi_8g_rx_pcs_dataout[38]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [38];
assign \w_hssi_8g_rx_pcs_dataout[39]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [39];
assign \w_hssi_8g_rx_pcs_dataout[40]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [40];
assign \w_hssi_8g_rx_pcs_dataout[41]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [41];
assign \w_hssi_8g_rx_pcs_dataout[42]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [42];
assign \w_hssi_8g_rx_pcs_dataout[43]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [43];
assign \w_hssi_8g_rx_pcs_dataout[44]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [44];
assign \w_hssi_8g_rx_pcs_dataout[45]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [45];
assign \w_hssi_8g_rx_pcs_dataout[46]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [46];
assign \w_hssi_8g_rx_pcs_dataout[47]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [47];
assign \w_hssi_8g_rx_pcs_dataout[48]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [48];
assign \w_hssi_8g_rx_pcs_dataout[49]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [49];
assign \w_hssi_8g_rx_pcs_dataout[50]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [50];
assign \w_hssi_8g_rx_pcs_dataout[51]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [51];
assign \w_hssi_8g_rx_pcs_dataout[52]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [52];
assign \w_hssi_8g_rx_pcs_dataout[53]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [53];
assign \w_hssi_8g_rx_pcs_dataout[54]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [54];
assign \w_hssi_8g_rx_pcs_dataout[55]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [55];
assign \w_hssi_8g_rx_pcs_dataout[56]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [56];
assign \w_hssi_8g_rx_pcs_dataout[57]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [57];
assign \w_hssi_8g_rx_pcs_dataout[58]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [58];
assign \w_hssi_8g_rx_pcs_dataout[59]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [59];
assign \w_hssi_8g_rx_pcs_dataout[60]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [60];
assign \w_hssi_8g_rx_pcs_dataout[61]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [61];
assign \w_hssi_8g_rx_pcs_dataout[62]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [62];
assign \w_hssi_8g_rx_pcs_dataout[63]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus [63];

assign \w_hssi_8g_rx_pcs_a1a2k1k2flag[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus [0];
assign \w_hssi_8g_rx_pcs_a1a2k1k2flag[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus [1];
assign \w_hssi_8g_rx_pcs_a1a2k1k2flag[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus [2];
assign \w_hssi_8g_rx_pcs_a1a2k1k2flag[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus [3];

assign \w_hssi_8g_rx_pcs_rxstatus[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RXSTATUS_bus [0];
assign \w_hssi_8g_rx_pcs_rxstatus[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RXSTATUS_bus [1];
assign \w_hssi_8g_rx_pcs_rxstatus[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RXSTATUS_bus [2];

assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [0];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [1];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [2];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [3];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [4];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [5];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [6];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [7];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [8];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [9];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [10];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [11];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [12];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [13];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [14];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [15];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [16];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [17];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [18];
assign \w_hssi_8g_rx_pcs_chnl_test_bus_out[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus [19];

assign \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_EIOS_DET_CDR_CTRL_bus [0];
assign \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_EIOS_DET_CDR_CTRL_bus [1];
assign \w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_EIOS_DET_CDR_CTRL_bus [2];

assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [7];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [8];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [9];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [10];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [11];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [12];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [13];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [14];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [15];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [16];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [17];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [18];
assign \w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus [19];

assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [7];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [8];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [9];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [10];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [11];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [12];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [13];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [14];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [15];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [16];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [17];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [18];
assign \w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus [19];

assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus [7];

assign \w_hssi_8g_rx_pcs_rx_blk_start[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus [0];
assign \w_hssi_8g_rx_pcs_rx_blk_start[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus [1];
assign \w_hssi_8g_rx_pcs_rx_blk_start[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus [2];
assign \w_hssi_8g_rx_pcs_rx_blk_start[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus [3];

assign \w_hssi_8g_rx_pcs_rx_sync_hdr[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_SYNC_HDR_bus [0];
assign \w_hssi_8g_rx_pcs_rx_sync_hdr[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_SYNC_HDR_bus [1];

assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [7];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [8];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [9];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [10];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [11];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [12];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [13];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [14];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [15];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [16];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [17];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [18];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [19];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [20];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [21];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [22];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [23];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [24];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [25];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [26];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [27];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [28];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [29];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [30];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [31];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [32];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [33];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [34];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [35];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [36];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [37];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [38];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [39];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [40];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [41];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [42];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [43];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [44];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [45];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [46];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [47];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [48];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [49];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [50];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [51];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [52];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [53];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [54];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [55];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [56];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [57];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [58];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [59];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [60];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [61];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [62];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [63];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [64];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [65];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [66];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [67];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [68];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [69];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [70];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [71];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [72];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [73];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [74];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [75];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [76];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [77];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [78];
assign \w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus [79];

assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [7];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [8];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [9];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [10];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [11];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [12];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [13];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [14];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [15];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [16];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [17];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [18];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [19];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [20];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [21];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [22];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [23];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [24];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [25];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [26];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [27];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [28];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [29];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [30];
assign \w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus [31];

assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus [7];

assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [0];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [1];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [2];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [3];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [4];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [5];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [6];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [7];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [8];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [9];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [10];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [11];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [12];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [13];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [14];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [15];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [16];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [17];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [18];
assign \w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19]  = \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus [19];

assign out_avmmreaddata_hssi_pipe_gen1_2[0] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_pipe_gen1_2[1] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_pipe_gen1_2[2] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_pipe_gen1_2[3] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_pipe_gen1_2[4] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_pipe_gen1_2[5] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_pipe_gen1_2[6] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_pipe_gen1_2[7] = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus [7];

assign \w_hssi_pipe_gen1_2_rxstatus[0]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_RXSTATUS_bus [0];
assign \w_hssi_pipe_gen1_2_rxstatus[1]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_RXSTATUS_bus [1];
assign \w_hssi_pipe_gen1_2_rxstatus[2]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_RXSTATUS_bus [2];

assign \w_hssi_pipe_gen1_2_current_coeff[0]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [0];
assign \w_hssi_pipe_gen1_2_current_coeff[1]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [1];
assign \w_hssi_pipe_gen1_2_current_coeff[2]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [2];
assign \w_hssi_pipe_gen1_2_current_coeff[3]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [3];
assign \w_hssi_pipe_gen1_2_current_coeff[4]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [4];
assign \w_hssi_pipe_gen1_2_current_coeff[5]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [5];
assign \w_hssi_pipe_gen1_2_current_coeff[6]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [6];
assign \w_hssi_pipe_gen1_2_current_coeff[7]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [7];
assign \w_hssi_pipe_gen1_2_current_coeff[8]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [8];
assign \w_hssi_pipe_gen1_2_current_coeff[9]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [9];
assign \w_hssi_pipe_gen1_2_current_coeff[10]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [10];
assign \w_hssi_pipe_gen1_2_current_coeff[11]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [11];
assign \w_hssi_pipe_gen1_2_current_coeff[12]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [12];
assign \w_hssi_pipe_gen1_2_current_coeff[13]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [13];
assign \w_hssi_pipe_gen1_2_current_coeff[14]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [14];
assign \w_hssi_pipe_gen1_2_current_coeff[15]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [15];
assign \w_hssi_pipe_gen1_2_current_coeff[16]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [16];
assign \w_hssi_pipe_gen1_2_current_coeff[17]  = \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus [17];

assign out_avmmreaddata_hssi_krfec_rx_pcs[0] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_krfec_rx_pcs[1] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_krfec_rx_pcs[2] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_krfec_rx_pcs[3] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_krfec_rx_pcs[4] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_krfec_rx_pcs[5] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_krfec_rx_pcs[6] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_krfec_rx_pcs[7] = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_krfec_rx_pcs_rx_control_out[0]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [0];
assign \w_hssi_krfec_rx_pcs_rx_control_out[1]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [1];
assign \w_hssi_krfec_rx_pcs_rx_control_out[2]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [2];
assign \w_hssi_krfec_rx_pcs_rx_control_out[3]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [3];
assign \w_hssi_krfec_rx_pcs_rx_control_out[4]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [4];
assign \w_hssi_krfec_rx_pcs_rx_control_out[5]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [5];
assign \w_hssi_krfec_rx_pcs_rx_control_out[6]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [6];
assign \w_hssi_krfec_rx_pcs_rx_control_out[7]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [7];
assign \w_hssi_krfec_rx_pcs_rx_control_out[8]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [8];
assign \w_hssi_krfec_rx_pcs_rx_control_out[9]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus [9];

assign \w_hssi_krfec_rx_pcs_rx_data_out[0]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [0];
assign \w_hssi_krfec_rx_pcs_rx_data_out[1]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [1];
assign \w_hssi_krfec_rx_pcs_rx_data_out[2]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [2];
assign \w_hssi_krfec_rx_pcs_rx_data_out[3]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [3];
assign \w_hssi_krfec_rx_pcs_rx_data_out[4]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [4];
assign \w_hssi_krfec_rx_pcs_rx_data_out[5]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [5];
assign \w_hssi_krfec_rx_pcs_rx_data_out[6]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [6];
assign \w_hssi_krfec_rx_pcs_rx_data_out[7]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [7];
assign \w_hssi_krfec_rx_pcs_rx_data_out[8]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [8];
assign \w_hssi_krfec_rx_pcs_rx_data_out[9]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [9];
assign \w_hssi_krfec_rx_pcs_rx_data_out[10]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [10];
assign \w_hssi_krfec_rx_pcs_rx_data_out[11]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [11];
assign \w_hssi_krfec_rx_pcs_rx_data_out[12]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [12];
assign \w_hssi_krfec_rx_pcs_rx_data_out[13]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [13];
assign \w_hssi_krfec_rx_pcs_rx_data_out[14]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [14];
assign \w_hssi_krfec_rx_pcs_rx_data_out[15]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [15];
assign \w_hssi_krfec_rx_pcs_rx_data_out[16]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [16];
assign \w_hssi_krfec_rx_pcs_rx_data_out[17]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [17];
assign \w_hssi_krfec_rx_pcs_rx_data_out[18]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [18];
assign \w_hssi_krfec_rx_pcs_rx_data_out[19]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [19];
assign \w_hssi_krfec_rx_pcs_rx_data_out[20]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [20];
assign \w_hssi_krfec_rx_pcs_rx_data_out[21]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [21];
assign \w_hssi_krfec_rx_pcs_rx_data_out[22]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [22];
assign \w_hssi_krfec_rx_pcs_rx_data_out[23]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [23];
assign \w_hssi_krfec_rx_pcs_rx_data_out[24]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [24];
assign \w_hssi_krfec_rx_pcs_rx_data_out[25]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [25];
assign \w_hssi_krfec_rx_pcs_rx_data_out[26]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [26];
assign \w_hssi_krfec_rx_pcs_rx_data_out[27]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [27];
assign \w_hssi_krfec_rx_pcs_rx_data_out[28]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [28];
assign \w_hssi_krfec_rx_pcs_rx_data_out[29]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [29];
assign \w_hssi_krfec_rx_pcs_rx_data_out[30]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [30];
assign \w_hssi_krfec_rx_pcs_rx_data_out[31]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [31];
assign \w_hssi_krfec_rx_pcs_rx_data_out[32]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [32];
assign \w_hssi_krfec_rx_pcs_rx_data_out[33]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [33];
assign \w_hssi_krfec_rx_pcs_rx_data_out[34]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [34];
assign \w_hssi_krfec_rx_pcs_rx_data_out[35]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [35];
assign \w_hssi_krfec_rx_pcs_rx_data_out[36]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [36];
assign \w_hssi_krfec_rx_pcs_rx_data_out[37]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [37];
assign \w_hssi_krfec_rx_pcs_rx_data_out[38]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [38];
assign \w_hssi_krfec_rx_pcs_rx_data_out[39]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [39];
assign \w_hssi_krfec_rx_pcs_rx_data_out[40]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [40];
assign \w_hssi_krfec_rx_pcs_rx_data_out[41]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [41];
assign \w_hssi_krfec_rx_pcs_rx_data_out[42]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [42];
assign \w_hssi_krfec_rx_pcs_rx_data_out[43]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [43];
assign \w_hssi_krfec_rx_pcs_rx_data_out[44]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [44];
assign \w_hssi_krfec_rx_pcs_rx_data_out[45]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [45];
assign \w_hssi_krfec_rx_pcs_rx_data_out[46]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [46];
assign \w_hssi_krfec_rx_pcs_rx_data_out[47]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [47];
assign \w_hssi_krfec_rx_pcs_rx_data_out[48]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [48];
assign \w_hssi_krfec_rx_pcs_rx_data_out[49]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [49];
assign \w_hssi_krfec_rx_pcs_rx_data_out[50]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [50];
assign \w_hssi_krfec_rx_pcs_rx_data_out[51]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [51];
assign \w_hssi_krfec_rx_pcs_rx_data_out[52]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [52];
assign \w_hssi_krfec_rx_pcs_rx_data_out[53]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [53];
assign \w_hssi_krfec_rx_pcs_rx_data_out[54]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [54];
assign \w_hssi_krfec_rx_pcs_rx_data_out[55]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [55];
assign \w_hssi_krfec_rx_pcs_rx_data_out[56]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [56];
assign \w_hssi_krfec_rx_pcs_rx_data_out[57]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [57];
assign \w_hssi_krfec_rx_pcs_rx_data_out[58]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [58];
assign \w_hssi_krfec_rx_pcs_rx_data_out[59]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [59];
assign \w_hssi_krfec_rx_pcs_rx_data_out[60]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [60];
assign \w_hssi_krfec_rx_pcs_rx_data_out[61]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [61];
assign \w_hssi_krfec_rx_pcs_rx_data_out[62]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [62];
assign \w_hssi_krfec_rx_pcs_rx_data_out[63]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus [63];

assign \w_hssi_krfec_rx_pcs_rx_data_status[0]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_STATUS_bus [0];
assign \w_hssi_krfec_rx_pcs_rx_data_status[1]  = \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_STATUS_bus [1];

assign out_avmmreaddata_hssi_rx_pcs_pma_interface[0] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[1] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[2] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[3] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[4] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[5] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[6] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_rx_pcs_pma_interface[7] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus [7];

assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [0];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [1];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [2];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [3];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [4];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [5];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [6];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [7];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [8];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [9];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [10];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [11];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [12];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [13];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [14];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [15];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [16];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [17];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [18];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [19];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [20];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [21];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [22];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [23];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [24];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [25];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [26];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [27];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [28];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [29];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [30];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [31];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [32];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [33];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [34];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [35];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [36];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [37];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [38];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [39];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [40];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [41];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [42];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [43];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [44];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [45];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [46];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [47];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [48];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [49];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [50];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [51];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [52];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [53];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [54];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [55];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [56];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [57];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [58];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [59];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [60];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [61];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [62];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus [63];

assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [0];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [1];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [2];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [3];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [4];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [5];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [6];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [7];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [8];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [9];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [10];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [11];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [12];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [13];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [14];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [15];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [16];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [17];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [18];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus [19];

assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [0];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [1];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [2];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [3];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [4];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [5];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [6];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [7];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [8];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [9];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [10];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [11];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [12];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [13];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [14];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [15];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [16];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [17];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [18];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [19];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [20];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [21];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [22];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [23];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [24];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [25];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [26];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [27];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [28];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [29];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [30];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus [31];

assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [0];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [1];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [2];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [3];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [4];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [5];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [6];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [7];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [8];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [9];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [10];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [11];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [12];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [13];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [14];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [15];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [16];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [17];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [18];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [19];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [20];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [21];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [22];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [23];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [24];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [25];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [26];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [27];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [28];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [29];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [30];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [31];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [32];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [33];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [34];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [35];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [36];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [37];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [38];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [39];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [40];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [41];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [42];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [43];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [44];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [45];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [46];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [47];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [48];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [49];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [50];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [51];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [52];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [53];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [54];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [55];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [56];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [57];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [58];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [59];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [60];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [61];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [62];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus [63];

assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [0];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [1];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [2];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [3];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [4];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [5];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [6];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [7];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [8];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [9];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [10];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [11];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [12];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [13];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [14];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [15];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [16];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [17];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [18];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [19];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [20];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [21];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [22];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [23];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [24];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [25];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [26];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [27];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [28];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [29];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [30];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [31];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [32];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [33];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [34];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [35];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [36];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [37];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [38];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [39];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [40];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [41];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [42];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [43];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [44];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [45];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [46];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [47];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [48];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [49];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [50];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [51];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [52];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [53];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [54];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [55];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [56];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [57];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [58];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [59];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [60];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [61];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [62];
assign \w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus [63];

assign out_pma_eye_monitor[0] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [0];
assign out_pma_eye_monitor[1] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [1];
assign out_pma_eye_monitor[2] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [2];
assign out_pma_eye_monitor[3] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [3];
assign out_pma_eye_monitor[4] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [4];
assign out_pma_eye_monitor[5] = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus [5];

assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [0];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [1];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [2];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [3];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [4];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [5];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [6];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [7];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [8];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [9];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [10];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [11];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [12];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [13];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [14];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [15];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [16];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [17];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [18];
assign \w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus [19];

assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [0];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [1];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [2];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [3];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [4];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [5];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [6];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [7];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [8];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [9];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [10];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [11];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [12];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [13];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [14];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [15];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [16];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [17];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [18];
assign \w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19]  = \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus [19];

assign out_avmmreaddata_hssi_8g_tx_pcs[0] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_8g_tx_pcs[1] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_8g_tx_pcs[2] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_8g_tx_pcs[3] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_8g_tx_pcs[4] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_8g_tx_pcs[5] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_8g_tx_pcs[6] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_8g_tx_pcs[7] = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_8g_tx_pcs_dataout[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [0];
assign \w_hssi_8g_tx_pcs_dataout[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [1];
assign \w_hssi_8g_tx_pcs_dataout[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [2];
assign \w_hssi_8g_tx_pcs_dataout[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [3];
assign \w_hssi_8g_tx_pcs_dataout[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [4];
assign \w_hssi_8g_tx_pcs_dataout[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [5];
assign \w_hssi_8g_tx_pcs_dataout[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [6];
assign \w_hssi_8g_tx_pcs_dataout[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [7];
assign \w_hssi_8g_tx_pcs_dataout[8]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [8];
assign \w_hssi_8g_tx_pcs_dataout[9]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [9];
assign \w_hssi_8g_tx_pcs_dataout[10]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [10];
assign \w_hssi_8g_tx_pcs_dataout[11]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [11];
assign \w_hssi_8g_tx_pcs_dataout[12]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [12];
assign \w_hssi_8g_tx_pcs_dataout[13]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [13];
assign \w_hssi_8g_tx_pcs_dataout[14]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [14];
assign \w_hssi_8g_tx_pcs_dataout[15]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [15];
assign \w_hssi_8g_tx_pcs_dataout[16]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [16];
assign \w_hssi_8g_tx_pcs_dataout[17]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [17];
assign \w_hssi_8g_tx_pcs_dataout[18]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [18];
assign \w_hssi_8g_tx_pcs_dataout[19]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus [19];

assign \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_NON_GRAY_EIDLEINFERSEL_bus [0];
assign \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_NON_GRAY_EIDLEINFERSEL_bus [1];
assign \w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_NON_GRAY_EIDLEINFERSEL_bus [2];

assign \w_hssi_8g_tx_pcs_phfifo_txmargin[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PHFIFO_TXMARGIN_bus [0];
assign \w_hssi_8g_tx_pcs_phfifo_txmargin[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PHFIFO_TXMARGIN_bus [1];
assign \w_hssi_8g_tx_pcs_phfifo_txmargin[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PHFIFO_TXMARGIN_bus [2];

assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [0];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [1];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [2];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [3];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [4];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [5];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [6];
assign \w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus [7];

assign \w_hssi_8g_tx_pcs_tx_blk_start_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_BLK_START_OUT_bus [0];

assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [0];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [1];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [2];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [3];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [4];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [5];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [6];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [7];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [8];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [9];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [10];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [11];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [12];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [13];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [14];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [15];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [16];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [17];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [18];
assign \w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus [19];

assign \w_hssi_8g_tx_pcs_tx_data_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [0];
assign \w_hssi_8g_tx_pcs_tx_data_out[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [1];
assign \w_hssi_8g_tx_pcs_tx_data_out[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [2];
assign \w_hssi_8g_tx_pcs_tx_data_out[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [3];
assign \w_hssi_8g_tx_pcs_tx_data_out[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [4];
assign \w_hssi_8g_tx_pcs_tx_data_out[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [5];
assign \w_hssi_8g_tx_pcs_tx_data_out[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [6];
assign \w_hssi_8g_tx_pcs_tx_data_out[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [7];
assign \w_hssi_8g_tx_pcs_tx_data_out[8]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [8];
assign \w_hssi_8g_tx_pcs_tx_data_out[9]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [9];
assign \w_hssi_8g_tx_pcs_tx_data_out[10]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [10];
assign \w_hssi_8g_tx_pcs_tx_data_out[11]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [11];
assign \w_hssi_8g_tx_pcs_tx_data_out[12]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [12];
assign \w_hssi_8g_tx_pcs_tx_data_out[13]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [13];
assign \w_hssi_8g_tx_pcs_tx_data_out[14]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [14];
assign \w_hssi_8g_tx_pcs_tx_data_out[15]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [15];
assign \w_hssi_8g_tx_pcs_tx_data_out[16]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [16];
assign \w_hssi_8g_tx_pcs_tx_data_out[17]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [17];
assign \w_hssi_8g_tx_pcs_tx_data_out[18]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [18];
assign \w_hssi_8g_tx_pcs_tx_data_out[19]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [19];
assign \w_hssi_8g_tx_pcs_tx_data_out[20]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [20];
assign \w_hssi_8g_tx_pcs_tx_data_out[21]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [21];
assign \w_hssi_8g_tx_pcs_tx_data_out[22]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [22];
assign \w_hssi_8g_tx_pcs_tx_data_out[23]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [23];
assign \w_hssi_8g_tx_pcs_tx_data_out[24]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [24];
assign \w_hssi_8g_tx_pcs_tx_data_out[25]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [25];
assign \w_hssi_8g_tx_pcs_tx_data_out[26]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [26];
assign \w_hssi_8g_tx_pcs_tx_data_out[27]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [27];
assign \w_hssi_8g_tx_pcs_tx_data_out[28]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [28];
assign \w_hssi_8g_tx_pcs_tx_data_out[29]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [29];
assign \w_hssi_8g_tx_pcs_tx_data_out[30]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [30];
assign \w_hssi_8g_tx_pcs_tx_data_out[31]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus [31];

assign \w_hssi_8g_tx_pcs_tx_data_valid_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_VALID_OUT_bus [0];

assign \w_hssi_8g_tx_pcs_tx_datak_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus [0];
assign \w_hssi_8g_tx_pcs_tx_datak_out[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus [1];
assign \w_hssi_8g_tx_pcs_tx_datak_out[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus [2];
assign \w_hssi_8g_tx_pcs_tx_datak_out[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus [3];

assign \w_hssi_8g_tx_pcs_tx_div_sync[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DIV_SYNC_bus [0];
assign \w_hssi_8g_tx_pcs_tx_div_sync[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DIV_SYNC_bus [1];

assign \w_hssi_8g_tx_pcs_tx_sync_hdr_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_SYNC_HDR_OUT_bus [0];
assign \w_hssi_8g_tx_pcs_tx_sync_hdr_out[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_SYNC_HDR_OUT_bus [1];

assign \w_hssi_8g_tx_pcs_tx_testbus[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [0];
assign \w_hssi_8g_tx_pcs_tx_testbus[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [1];
assign \w_hssi_8g_tx_pcs_tx_testbus[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [2];
assign \w_hssi_8g_tx_pcs_tx_testbus[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [3];
assign \w_hssi_8g_tx_pcs_tx_testbus[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [4];
assign \w_hssi_8g_tx_pcs_tx_testbus[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [5];
assign \w_hssi_8g_tx_pcs_tx_testbus[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [6];
assign \w_hssi_8g_tx_pcs_tx_testbus[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [7];
assign \w_hssi_8g_tx_pcs_tx_testbus[8]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [8];
assign \w_hssi_8g_tx_pcs_tx_testbus[9]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [9];
assign \w_hssi_8g_tx_pcs_tx_testbus[10]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [10];
assign \w_hssi_8g_tx_pcs_tx_testbus[11]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [11];
assign \w_hssi_8g_tx_pcs_tx_testbus[12]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [12];
assign \w_hssi_8g_tx_pcs_tx_testbus[13]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [13];
assign \w_hssi_8g_tx_pcs_tx_testbus[14]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [14];
assign \w_hssi_8g_tx_pcs_tx_testbus[15]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [15];
assign \w_hssi_8g_tx_pcs_tx_testbus[16]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [16];
assign \w_hssi_8g_tx_pcs_tx_testbus[17]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [17];
assign \w_hssi_8g_tx_pcs_tx_testbus[18]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [18];
assign \w_hssi_8g_tx_pcs_tx_testbus[19]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus [19];

assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [0];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [1];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [2];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [3];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [4];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [5];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [6];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [7];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [8];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [9];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [10];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [11];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [12];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [13];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [14];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [15];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [16];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [17];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [18];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [19];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [20];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [21];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [22];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [23];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [24];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [25];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [26];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [27];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [28];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [29];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [30];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [31];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [32];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [33];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [34];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [35];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [36];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [37];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [38];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [39];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [40];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [41];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [42];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [43];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [44];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [45];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [46];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [47];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [48];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [49];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [50];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [51];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [52];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [53];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [54];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [55];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [56];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [57];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [58];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [59];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [60];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [61];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [62];
assign \w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus [63];

assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [0];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [1];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [2];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [3];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [4];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [5];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [6];
assign \w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus [7];

assign \w_hssi_8g_tx_pcs_pipe_power_down_out[0]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PIPE_POWER_DOWN_OUT_bus [0];
assign \w_hssi_8g_tx_pcs_pipe_power_down_out[1]  = \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PIPE_POWER_DOWN_OUT_bus [1];

assign \w_hssi_10g_tx_pcs_tx_pma_data[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [0];
assign \w_hssi_10g_tx_pcs_tx_pma_data[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [1];
assign \w_hssi_10g_tx_pcs_tx_pma_data[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [2];
assign \w_hssi_10g_tx_pcs_tx_pma_data[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [3];
assign \w_hssi_10g_tx_pcs_tx_pma_data[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [4];
assign \w_hssi_10g_tx_pcs_tx_pma_data[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [5];
assign \w_hssi_10g_tx_pcs_tx_pma_data[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [6];
assign \w_hssi_10g_tx_pcs_tx_pma_data[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [7];
assign \w_hssi_10g_tx_pcs_tx_pma_data[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [8];
assign \w_hssi_10g_tx_pcs_tx_pma_data[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [9];
assign \w_hssi_10g_tx_pcs_tx_pma_data[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [10];
assign \w_hssi_10g_tx_pcs_tx_pma_data[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [11];
assign \w_hssi_10g_tx_pcs_tx_pma_data[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [12];
assign \w_hssi_10g_tx_pcs_tx_pma_data[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [13];
assign \w_hssi_10g_tx_pcs_tx_pma_data[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [14];
assign \w_hssi_10g_tx_pcs_tx_pma_data[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [15];
assign \w_hssi_10g_tx_pcs_tx_pma_data[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [16];
assign \w_hssi_10g_tx_pcs_tx_pma_data[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [17];
assign \w_hssi_10g_tx_pcs_tx_pma_data[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [18];
assign \w_hssi_10g_tx_pcs_tx_pma_data[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [19];
assign \w_hssi_10g_tx_pcs_tx_pma_data[20]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [20];
assign \w_hssi_10g_tx_pcs_tx_pma_data[21]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [21];
assign \w_hssi_10g_tx_pcs_tx_pma_data[22]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [22];
assign \w_hssi_10g_tx_pcs_tx_pma_data[23]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [23];
assign \w_hssi_10g_tx_pcs_tx_pma_data[24]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [24];
assign \w_hssi_10g_tx_pcs_tx_pma_data[25]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [25];
assign \w_hssi_10g_tx_pcs_tx_pma_data[26]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [26];
assign \w_hssi_10g_tx_pcs_tx_pma_data[27]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [27];
assign \w_hssi_10g_tx_pcs_tx_pma_data[28]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [28];
assign \w_hssi_10g_tx_pcs_tx_pma_data[29]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [29];
assign \w_hssi_10g_tx_pcs_tx_pma_data[30]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [30];
assign \w_hssi_10g_tx_pcs_tx_pma_data[31]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [31];
assign \w_hssi_10g_tx_pcs_tx_pma_data[32]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [32];
assign \w_hssi_10g_tx_pcs_tx_pma_data[33]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [33];
assign \w_hssi_10g_tx_pcs_tx_pma_data[34]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [34];
assign \w_hssi_10g_tx_pcs_tx_pma_data[35]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [35];
assign \w_hssi_10g_tx_pcs_tx_pma_data[36]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [36];
assign \w_hssi_10g_tx_pcs_tx_pma_data[37]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [37];
assign \w_hssi_10g_tx_pcs_tx_pma_data[38]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [38];
assign \w_hssi_10g_tx_pcs_tx_pma_data[39]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [39];
assign \w_hssi_10g_tx_pcs_tx_pma_data[40]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [40];
assign \w_hssi_10g_tx_pcs_tx_pma_data[41]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [41];
assign \w_hssi_10g_tx_pcs_tx_pma_data[42]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [42];
assign \w_hssi_10g_tx_pcs_tx_pma_data[43]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [43];
assign \w_hssi_10g_tx_pcs_tx_pma_data[44]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [44];
assign \w_hssi_10g_tx_pcs_tx_pma_data[45]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [45];
assign \w_hssi_10g_tx_pcs_tx_pma_data[46]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [46];
assign \w_hssi_10g_tx_pcs_tx_pma_data[47]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [47];
assign \w_hssi_10g_tx_pcs_tx_pma_data[48]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [48];
assign \w_hssi_10g_tx_pcs_tx_pma_data[49]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [49];
assign \w_hssi_10g_tx_pcs_tx_pma_data[50]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [50];
assign \w_hssi_10g_tx_pcs_tx_pma_data[51]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [51];
assign \w_hssi_10g_tx_pcs_tx_pma_data[52]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [52];
assign \w_hssi_10g_tx_pcs_tx_pma_data[53]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [53];
assign \w_hssi_10g_tx_pcs_tx_pma_data[54]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [54];
assign \w_hssi_10g_tx_pcs_tx_pma_data[55]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [55];
assign \w_hssi_10g_tx_pcs_tx_pma_data[56]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [56];
assign \w_hssi_10g_tx_pcs_tx_pma_data[57]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [57];
assign \w_hssi_10g_tx_pcs_tx_pma_data[58]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [58];
assign \w_hssi_10g_tx_pcs_tx_pma_data[59]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [59];
assign \w_hssi_10g_tx_pcs_tx_pma_data[60]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [60];
assign \w_hssi_10g_tx_pcs_tx_pma_data[61]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [61];
assign \w_hssi_10g_tx_pcs_tx_pma_data[62]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [62];
assign \w_hssi_10g_tx_pcs_tx_pma_data[63]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus [63];

assign out_avmmreaddata_hssi_10g_tx_pcs[0] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_10g_tx_pcs[1] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_10g_tx_pcs[2] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_10g_tx_pcs[3] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_10g_tx_pcs[4] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_10g_tx_pcs[5] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_10g_tx_pcs[6] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_10g_tx_pcs[7] = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [0];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [1];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [2];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [3];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [4];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [5];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [6];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [7];
assign \w_hssi_10g_tx_pcs_tx_control_out_krfec[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus [8];

assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [0];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [1];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [2];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [3];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [4];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [5];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [6];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [7];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [8];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [9];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [10];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [11];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [12];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [13];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [14];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [15];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [16];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [17];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [18];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [19];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[20]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [20];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[21]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [21];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[22]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [22];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[23]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [23];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[24]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [24];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[25]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [25];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[26]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [26];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[27]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [27];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[28]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [28];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[29]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [29];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[30]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [30];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[31]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [31];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[32]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [32];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[33]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [33];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[34]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [34];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[35]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [35];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[36]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [36];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[37]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [37];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[38]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [38];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[39]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [39];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[40]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [40];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[41]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [41];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[42]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [42];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[43]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [43];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[44]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [44];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[45]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [45];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[46]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [46];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[47]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [47];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[48]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [48];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[49]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [49];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[50]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [50];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[51]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [51];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[52]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [52];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[53]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [53];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[54]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [54];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[55]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [55];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[56]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [56];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[57]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [57];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[58]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [58];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[59]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [59];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[60]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [60];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[61]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [61];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[62]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [62];
assign \w_hssi_10g_tx_pcs_tx_data_out_krfec[63]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus [63];

assign \w_hssi_10g_tx_pcs_tx_fifo_num[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus [0];
assign \w_hssi_10g_tx_pcs_tx_fifo_num[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus [1];
assign \w_hssi_10g_tx_pcs_tx_fifo_num[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus [2];
assign \w_hssi_10g_tx_pcs_tx_fifo_num[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus [3];

assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [0];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [1];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [2];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [3];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [4];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [5];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [6];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [7];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [8];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [9];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [10];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [11];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [12];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [13];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [14];
assign \w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus [15];

assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [0];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [1];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [2];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [3];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [4];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [5];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [6];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [7];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [8];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [9];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [10];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [11];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [12];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [13];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [14];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [15];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [16];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [17];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [18];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [19];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[20]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [20];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[21]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [21];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[22]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [22];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[23]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [23];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[24]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [24];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[25]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [25];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[26]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [26];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[27]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [27];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[28]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [28];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[29]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [29];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[30]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [30];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[31]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [31];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[32]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [32];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[33]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [33];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[34]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [34];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[35]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [35];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[36]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [36];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[37]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [37];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[38]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [38];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[39]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [39];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[40]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [40];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[41]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [41];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[42]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [42];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[43]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [43];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[44]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [44];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[45]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [45];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[46]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [46];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[47]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [47];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[48]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [48];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[49]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [49];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[50]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [50];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[51]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [51];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[52]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [52];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[53]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [53];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[54]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [54];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[55]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [55];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[56]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [56];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[57]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [57];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[58]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [58];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[59]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [59];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[60]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [60];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[61]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [61];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[62]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [62];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[63]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [63];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[64]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [64];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[65]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [65];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[66]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [66];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[67]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [67];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[68]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [68];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[69]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [69];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[70]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [70];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[71]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [71];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data[72]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus [72];

assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [0];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [1];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [2];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [3];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [4];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [5];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [6];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [7];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [8];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [9];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [10];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [11];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [12];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [13];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [14];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [15];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [16];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [17];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [18];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [19];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [20];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [21];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [22];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [23];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [24];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [25];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [26];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [27];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [28];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [29];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [30];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [31];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [32];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [33];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [34];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [35];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [36];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [37];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [38];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [39];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [40];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [41];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [42];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [43];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [44];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [45];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [46];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [47];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [48];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [49];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [50];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [51];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [52];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [53];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [54];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [55];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [56];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [57];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [58];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [59];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [60];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [61];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [62];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [63];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [64];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [65];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [66];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [67];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [68];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [69];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [70];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [71];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus [72];

assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [0];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [1];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [2];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [3];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [4];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [5];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [6];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [7];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [8];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [9];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [10];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [11];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [12];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [13];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [14];
assign \w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus [15];

assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [0];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [1];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [2];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [3];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [4];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [5];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [6];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [7];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [8];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [9];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [10];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [11];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [12];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [13];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [14];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [15];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [16];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [17];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [18];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [19];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[20]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [20];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[21]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [21];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[22]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [22];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[23]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [23];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[24]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [24];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[25]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [25];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[26]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [26];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[27]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [27];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[28]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [28];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[29]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [29];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[30]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [30];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[31]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [31];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[32]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [32];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[33]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [33];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[34]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [34];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[35]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [35];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[36]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [36];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[37]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [37];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[38]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [38];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[39]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [39];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[40]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [40];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[41]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [41];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[42]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [42];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[43]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [43];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[44]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [44];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[45]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [45];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[46]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [46];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[47]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [47];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[48]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [48];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[49]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [49];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[50]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [50];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[51]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [51];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[52]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [52];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[53]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [53];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[54]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [54];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[55]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [55];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[56]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [56];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[57]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [57];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[58]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [58];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[59]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [59];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[60]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [60];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[61]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [61];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[62]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [62];
assign \w_hssi_10g_tx_pcs_tx_pma_gating_val[63]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus [63];

assign \w_hssi_10g_tx_pcs_tx_test_data[0]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [0];
assign \w_hssi_10g_tx_pcs_tx_test_data[1]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [1];
assign \w_hssi_10g_tx_pcs_tx_test_data[2]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [2];
assign \w_hssi_10g_tx_pcs_tx_test_data[3]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [3];
assign \w_hssi_10g_tx_pcs_tx_test_data[4]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [4];
assign \w_hssi_10g_tx_pcs_tx_test_data[5]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [5];
assign \w_hssi_10g_tx_pcs_tx_test_data[6]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [6];
assign \w_hssi_10g_tx_pcs_tx_test_data[7]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [7];
assign \w_hssi_10g_tx_pcs_tx_test_data[8]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [8];
assign \w_hssi_10g_tx_pcs_tx_test_data[9]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [9];
assign \w_hssi_10g_tx_pcs_tx_test_data[10]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [10];
assign \w_hssi_10g_tx_pcs_tx_test_data[11]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [11];
assign \w_hssi_10g_tx_pcs_tx_test_data[12]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [12];
assign \w_hssi_10g_tx_pcs_tx_test_data[13]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [13];
assign \w_hssi_10g_tx_pcs_tx_test_data[14]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [14];
assign \w_hssi_10g_tx_pcs_tx_test_data[15]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [15];
assign \w_hssi_10g_tx_pcs_tx_test_data[16]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [16];
assign \w_hssi_10g_tx_pcs_tx_test_data[17]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [17];
assign \w_hssi_10g_tx_pcs_tx_test_data[18]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [18];
assign \w_hssi_10g_tx_pcs_tx_test_data[19]  = \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus [19];

assign \w_hssi_gen3_rx_pcs_data_out[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [0];
assign \w_hssi_gen3_rx_pcs_data_out[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [1];
assign \w_hssi_gen3_rx_pcs_data_out[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [2];
assign \w_hssi_gen3_rx_pcs_data_out[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [3];
assign \w_hssi_gen3_rx_pcs_data_out[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [4];
assign \w_hssi_gen3_rx_pcs_data_out[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [5];
assign \w_hssi_gen3_rx_pcs_data_out[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [6];
assign \w_hssi_gen3_rx_pcs_data_out[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [7];
assign \w_hssi_gen3_rx_pcs_data_out[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [8];
assign \w_hssi_gen3_rx_pcs_data_out[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [9];
assign \w_hssi_gen3_rx_pcs_data_out[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [10];
assign \w_hssi_gen3_rx_pcs_data_out[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [11];
assign \w_hssi_gen3_rx_pcs_data_out[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [12];
assign \w_hssi_gen3_rx_pcs_data_out[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [13];
assign \w_hssi_gen3_rx_pcs_data_out[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [14];
assign \w_hssi_gen3_rx_pcs_data_out[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [15];
assign \w_hssi_gen3_rx_pcs_data_out[16]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [16];
assign \w_hssi_gen3_rx_pcs_data_out[17]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [17];
assign \w_hssi_gen3_rx_pcs_data_out[18]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [18];
assign \w_hssi_gen3_rx_pcs_data_out[19]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [19];
assign \w_hssi_gen3_rx_pcs_data_out[20]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [20];
assign \w_hssi_gen3_rx_pcs_data_out[21]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [21];
assign \w_hssi_gen3_rx_pcs_data_out[22]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [22];
assign \w_hssi_gen3_rx_pcs_data_out[23]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [23];
assign \w_hssi_gen3_rx_pcs_data_out[24]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [24];
assign \w_hssi_gen3_rx_pcs_data_out[25]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [25];
assign \w_hssi_gen3_rx_pcs_data_out[26]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [26];
assign \w_hssi_gen3_rx_pcs_data_out[27]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [27];
assign \w_hssi_gen3_rx_pcs_data_out[28]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [28];
assign \w_hssi_gen3_rx_pcs_data_out[29]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [29];
assign \w_hssi_gen3_rx_pcs_data_out[30]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [30];
assign \w_hssi_gen3_rx_pcs_data_out[31]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus [31];

assign out_avmmreaddata_hssi_gen3_rx_pcs[0] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_gen3_rx_pcs[1] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_gen3_rx_pcs[2] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_gen3_rx_pcs[3] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_gen3_rx_pcs[4] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_gen3_rx_pcs[5] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_gen3_rx_pcs[6] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_gen3_rx_pcs[7] = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_gen3_rx_pcs_lpbk_data[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [0];
assign \w_hssi_gen3_rx_pcs_lpbk_data[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [1];
assign \w_hssi_gen3_rx_pcs_lpbk_data[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [2];
assign \w_hssi_gen3_rx_pcs_lpbk_data[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [3];
assign \w_hssi_gen3_rx_pcs_lpbk_data[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [4];
assign \w_hssi_gen3_rx_pcs_lpbk_data[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [5];
assign \w_hssi_gen3_rx_pcs_lpbk_data[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [6];
assign \w_hssi_gen3_rx_pcs_lpbk_data[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [7];
assign \w_hssi_gen3_rx_pcs_lpbk_data[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [8];
assign \w_hssi_gen3_rx_pcs_lpbk_data[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [9];
assign \w_hssi_gen3_rx_pcs_lpbk_data[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [10];
assign \w_hssi_gen3_rx_pcs_lpbk_data[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [11];
assign \w_hssi_gen3_rx_pcs_lpbk_data[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [12];
assign \w_hssi_gen3_rx_pcs_lpbk_data[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [13];
assign \w_hssi_gen3_rx_pcs_lpbk_data[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [14];
assign \w_hssi_gen3_rx_pcs_lpbk_data[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [15];
assign \w_hssi_gen3_rx_pcs_lpbk_data[16]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [16];
assign \w_hssi_gen3_rx_pcs_lpbk_data[17]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [17];
assign \w_hssi_gen3_rx_pcs_lpbk_data[18]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [18];
assign \w_hssi_gen3_rx_pcs_lpbk_data[19]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [19];
assign \w_hssi_gen3_rx_pcs_lpbk_data[20]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [20];
assign \w_hssi_gen3_rx_pcs_lpbk_data[21]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [21];
assign \w_hssi_gen3_rx_pcs_lpbk_data[22]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [22];
assign \w_hssi_gen3_rx_pcs_lpbk_data[23]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [23];
assign \w_hssi_gen3_rx_pcs_lpbk_data[24]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [24];
assign \w_hssi_gen3_rx_pcs_lpbk_data[25]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [25];
assign \w_hssi_gen3_rx_pcs_lpbk_data[26]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [26];
assign \w_hssi_gen3_rx_pcs_lpbk_data[27]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [27];
assign \w_hssi_gen3_rx_pcs_lpbk_data[28]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [28];
assign \w_hssi_gen3_rx_pcs_lpbk_data[29]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [29];
assign \w_hssi_gen3_rx_pcs_lpbk_data[30]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [30];
assign \w_hssi_gen3_rx_pcs_lpbk_data[31]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [31];
assign \w_hssi_gen3_rx_pcs_lpbk_data[32]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [32];
assign \w_hssi_gen3_rx_pcs_lpbk_data[33]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus [33];

assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [0];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [1];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [2];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [3];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [4];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [5];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [6];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [7];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [8];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [9];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [10];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [11];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [12];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [13];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [14];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus [15];

assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [0];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [1];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [2];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [3];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [4];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [5];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [6];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [7];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [8];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [9];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [10];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [11];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [12];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [13];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [14];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [15];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [16];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [17];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [18];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [19];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [20];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [21];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [22];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [23];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [24];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [25];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [26];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [27];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [28];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [29];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [30];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [31];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [32];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [33];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [34];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [35];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [36];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [37];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [38];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus [39];

assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [0];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [1];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [2];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [3];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [4];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [5];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [6];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [7];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [8];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [9];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [10];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [11];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [12];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [13];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [14];
assign \w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus [15];

assign \w_hssi_gen3_rx_pcs_rx_test_out[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [0];
assign \w_hssi_gen3_rx_pcs_rx_test_out[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [1];
assign \w_hssi_gen3_rx_pcs_rx_test_out[2]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [2];
assign \w_hssi_gen3_rx_pcs_rx_test_out[3]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [3];
assign \w_hssi_gen3_rx_pcs_rx_test_out[4]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [4];
assign \w_hssi_gen3_rx_pcs_rx_test_out[5]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [5];
assign \w_hssi_gen3_rx_pcs_rx_test_out[6]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [6];
assign \w_hssi_gen3_rx_pcs_rx_test_out[7]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [7];
assign \w_hssi_gen3_rx_pcs_rx_test_out[8]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [8];
assign \w_hssi_gen3_rx_pcs_rx_test_out[9]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [9];
assign \w_hssi_gen3_rx_pcs_rx_test_out[10]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [10];
assign \w_hssi_gen3_rx_pcs_rx_test_out[11]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [11];
assign \w_hssi_gen3_rx_pcs_rx_test_out[12]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [12];
assign \w_hssi_gen3_rx_pcs_rx_test_out[13]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [13];
assign \w_hssi_gen3_rx_pcs_rx_test_out[14]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [14];
assign \w_hssi_gen3_rx_pcs_rx_test_out[15]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [15];
assign \w_hssi_gen3_rx_pcs_rx_test_out[16]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [16];
assign \w_hssi_gen3_rx_pcs_rx_test_out[17]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [17];
assign \w_hssi_gen3_rx_pcs_rx_test_out[18]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [18];
assign \w_hssi_gen3_rx_pcs_rx_test_out[19]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus [19];

assign \w_hssi_gen3_rx_pcs_sync_hdr[0]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_SYNC_HDR_bus [0];
assign \w_hssi_gen3_rx_pcs_sync_hdr[1]  = \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_SYNC_HDR_bus [1];

assign \w_hssi_pipe_gen3_test_out[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [0];
assign \w_hssi_pipe_gen3_test_out[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [1];
assign \w_hssi_pipe_gen3_test_out[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [2];
assign \w_hssi_pipe_gen3_test_out[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [3];
assign \w_hssi_pipe_gen3_test_out[4]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [4];
assign \w_hssi_pipe_gen3_test_out[5]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [5];
assign \w_hssi_pipe_gen3_test_out[6]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [6];
assign \w_hssi_pipe_gen3_test_out[7]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [7];
assign \w_hssi_pipe_gen3_test_out[8]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [8];
assign \w_hssi_pipe_gen3_test_out[9]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [9];
assign \w_hssi_pipe_gen3_test_out[10]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [10];
assign \w_hssi_pipe_gen3_test_out[11]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [11];
assign \w_hssi_pipe_gen3_test_out[12]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [12];
assign \w_hssi_pipe_gen3_test_out[13]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [13];
assign \w_hssi_pipe_gen3_test_out[14]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [14];
assign \w_hssi_pipe_gen3_test_out[15]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [15];
assign \w_hssi_pipe_gen3_test_out[16]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [16];
assign \w_hssi_pipe_gen3_test_out[17]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [17];
assign \w_hssi_pipe_gen3_test_out[18]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [18];
assign \w_hssi_pipe_gen3_test_out[19]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus [19];

assign out_avmmreaddata_hssi_pipe_gen3[0] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_pipe_gen3[1] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_pipe_gen3[2] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_pipe_gen3[3] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_pipe_gen3[4] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_pipe_gen3[5] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_pipe_gen3[6] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_pipe_gen3[7] = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus [7];

assign \w_hssi_pipe_gen3_rxstatus[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXSTATUS_bus [0];
assign \w_hssi_pipe_gen3_rxstatus[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXSTATUS_bus [1];
assign \w_hssi_pipe_gen3_rxstatus[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXSTATUS_bus [2];

assign \w_hssi_pipe_gen3_rx_blk_start[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus [0];
assign \w_hssi_pipe_gen3_rx_blk_start[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus [1];
assign \w_hssi_pipe_gen3_rx_blk_start[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus [2];
assign \w_hssi_pipe_gen3_rx_blk_start[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus [3];

assign \w_hssi_pipe_gen3_rx_sync_hdr[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_SYNC_HDR_bus [0];
assign \w_hssi_pipe_gen3_rx_sync_hdr[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_SYNC_HDR_bus [1];

assign \w_hssi_pipe_gen3_pma_current_coeff[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [0];
assign \w_hssi_pipe_gen3_pma_current_coeff[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [1];
assign \w_hssi_pipe_gen3_pma_current_coeff[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [2];
assign \w_hssi_pipe_gen3_pma_current_coeff[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [3];
assign \w_hssi_pipe_gen3_pma_current_coeff[4]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [4];
assign \w_hssi_pipe_gen3_pma_current_coeff[5]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [5];
assign \w_hssi_pipe_gen3_pma_current_coeff[6]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [6];
assign \w_hssi_pipe_gen3_pma_current_coeff[7]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [7];
assign \w_hssi_pipe_gen3_pma_current_coeff[8]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [8];
assign \w_hssi_pipe_gen3_pma_current_coeff[9]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [9];
assign \w_hssi_pipe_gen3_pma_current_coeff[10]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [10];
assign \w_hssi_pipe_gen3_pma_current_coeff[11]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [11];
assign \w_hssi_pipe_gen3_pma_current_coeff[12]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [12];
assign \w_hssi_pipe_gen3_pma_current_coeff[13]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [13];
assign \w_hssi_pipe_gen3_pma_current_coeff[14]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [14];
assign \w_hssi_pipe_gen3_pma_current_coeff[15]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [15];
assign \w_hssi_pipe_gen3_pma_current_coeff[16]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [16];
assign \w_hssi_pipe_gen3_pma_current_coeff[17]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus [17];

assign \w_hssi_pipe_gen3_pma_current_rxpreset[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_RXPRESET_bus [0];
assign \w_hssi_pipe_gen3_pma_current_rxpreset[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_RXPRESET_bus [1];
assign \w_hssi_pipe_gen3_pma_current_rxpreset[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_RXPRESET_bus [2];

assign \w_hssi_pipe_gen3_rxd_8gpcs_out[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [0];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [1];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [2];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [3];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[4]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [4];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[5]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [5];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[6]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [6];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[7]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [7];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[8]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [8];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[9]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [9];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[10]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [10];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[11]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [11];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[12]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [12];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[13]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [13];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[14]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [14];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[15]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [15];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[16]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [16];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[17]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [17];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[18]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [18];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[19]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [19];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[20]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [20];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[21]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [21];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[22]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [22];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[23]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [23];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[24]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [24];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[25]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [25];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[26]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [26];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[27]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [27];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[28]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [28];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[29]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [29];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[30]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [30];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[31]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [31];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[32]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [32];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[33]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [33];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[34]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [34];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[35]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [35];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[36]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [36];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[37]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [37];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[38]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [38];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[39]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [39];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[40]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [40];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[41]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [41];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[42]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [42];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[43]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [43];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[44]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [44];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[45]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [45];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[46]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [46];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[47]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [47];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[48]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [48];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[49]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [49];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[50]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [50];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[51]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [51];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[52]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [52];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[53]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [53];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[54]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [54];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[55]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [55];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[56]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [56];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[57]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [57];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[58]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [58];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[59]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [59];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[60]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [60];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[61]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [61];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[62]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [62];
assign \w_hssi_pipe_gen3_rxd_8gpcs_out[63]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus [63];

assign \w_hssi_pipe_gen3_rxdataskip[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus [0];
assign \w_hssi_pipe_gen3_rxdataskip[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus [1];
assign \w_hssi_pipe_gen3_rxdataskip[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus [2];
assign \w_hssi_pipe_gen3_rxdataskip[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus [3];

assign \w_hssi_pipe_gen3_tx_sync_hdr_int[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TX_SYNC_HDR_INT_bus [0];
assign \w_hssi_pipe_gen3_tx_sync_hdr_int[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TX_SYNC_HDR_INT_bus [1];

assign \w_hssi_pipe_gen3_txdata_int[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [0];
assign \w_hssi_pipe_gen3_txdata_int[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [1];
assign \w_hssi_pipe_gen3_txdata_int[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [2];
assign \w_hssi_pipe_gen3_txdata_int[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [3];
assign \w_hssi_pipe_gen3_txdata_int[4]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [4];
assign \w_hssi_pipe_gen3_txdata_int[5]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [5];
assign \w_hssi_pipe_gen3_txdata_int[6]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [6];
assign \w_hssi_pipe_gen3_txdata_int[7]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [7];
assign \w_hssi_pipe_gen3_txdata_int[8]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [8];
assign \w_hssi_pipe_gen3_txdata_int[9]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [9];
assign \w_hssi_pipe_gen3_txdata_int[10]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [10];
assign \w_hssi_pipe_gen3_txdata_int[11]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [11];
assign \w_hssi_pipe_gen3_txdata_int[12]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [12];
assign \w_hssi_pipe_gen3_txdata_int[13]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [13];
assign \w_hssi_pipe_gen3_txdata_int[14]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [14];
assign \w_hssi_pipe_gen3_txdata_int[15]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [15];
assign \w_hssi_pipe_gen3_txdata_int[16]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [16];
assign \w_hssi_pipe_gen3_txdata_int[17]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [17];
assign \w_hssi_pipe_gen3_txdata_int[18]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [18];
assign \w_hssi_pipe_gen3_txdata_int[19]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [19];
assign \w_hssi_pipe_gen3_txdata_int[20]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [20];
assign \w_hssi_pipe_gen3_txdata_int[21]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [21];
assign \w_hssi_pipe_gen3_txdata_int[22]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [22];
assign \w_hssi_pipe_gen3_txdata_int[23]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [23];
assign \w_hssi_pipe_gen3_txdata_int[24]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [24];
assign \w_hssi_pipe_gen3_txdata_int[25]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [25];
assign \w_hssi_pipe_gen3_txdata_int[26]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [26];
assign \w_hssi_pipe_gen3_txdata_int[27]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [27];
assign \w_hssi_pipe_gen3_txdata_int[28]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [28];
assign \w_hssi_pipe_gen3_txdata_int[29]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [29];
assign \w_hssi_pipe_gen3_txdata_int[30]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [30];
assign \w_hssi_pipe_gen3_txdata_int[31]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus [31];

assign \w_hssi_pipe_gen3_txdatak_int[0]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus [0];
assign \w_hssi_pipe_gen3_txdatak_int[1]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus [1];
assign \w_hssi_pipe_gen3_txdatak_int[2]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus [2];
assign \w_hssi_pipe_gen3_txdatak_int[3]  = \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus [3];

assign \w_hssi_gen3_tx_pcs_data_out[0]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [0];
assign \w_hssi_gen3_tx_pcs_data_out[1]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [1];
assign \w_hssi_gen3_tx_pcs_data_out[2]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [2];
assign \w_hssi_gen3_tx_pcs_data_out[3]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [3];
assign \w_hssi_gen3_tx_pcs_data_out[4]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [4];
assign \w_hssi_gen3_tx_pcs_data_out[5]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [5];
assign \w_hssi_gen3_tx_pcs_data_out[6]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [6];
assign \w_hssi_gen3_tx_pcs_data_out[7]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [7];
assign \w_hssi_gen3_tx_pcs_data_out[8]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [8];
assign \w_hssi_gen3_tx_pcs_data_out[9]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [9];
assign \w_hssi_gen3_tx_pcs_data_out[10]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [10];
assign \w_hssi_gen3_tx_pcs_data_out[11]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [11];
assign \w_hssi_gen3_tx_pcs_data_out[12]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [12];
assign \w_hssi_gen3_tx_pcs_data_out[13]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [13];
assign \w_hssi_gen3_tx_pcs_data_out[14]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [14];
assign \w_hssi_gen3_tx_pcs_data_out[15]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [15];
assign \w_hssi_gen3_tx_pcs_data_out[16]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [16];
assign \w_hssi_gen3_tx_pcs_data_out[17]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [17];
assign \w_hssi_gen3_tx_pcs_data_out[18]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [18];
assign \w_hssi_gen3_tx_pcs_data_out[19]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [19];
assign \w_hssi_gen3_tx_pcs_data_out[20]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [20];
assign \w_hssi_gen3_tx_pcs_data_out[21]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [21];
assign \w_hssi_gen3_tx_pcs_data_out[22]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [22];
assign \w_hssi_gen3_tx_pcs_data_out[23]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [23];
assign \w_hssi_gen3_tx_pcs_data_out[24]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [24];
assign \w_hssi_gen3_tx_pcs_data_out[25]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [25];
assign \w_hssi_gen3_tx_pcs_data_out[26]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [26];
assign \w_hssi_gen3_tx_pcs_data_out[27]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [27];
assign \w_hssi_gen3_tx_pcs_data_out[28]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [28];
assign \w_hssi_gen3_tx_pcs_data_out[29]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [29];
assign \w_hssi_gen3_tx_pcs_data_out[30]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [30];
assign \w_hssi_gen3_tx_pcs_data_out[31]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus [31];

assign out_avmmreaddata_hssi_gen3_tx_pcs[0] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_gen3_tx_pcs[1] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_gen3_tx_pcs[2] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_gen3_tx_pcs[3] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_gen3_tx_pcs[4] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_gen3_tx_pcs[5] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_gen3_tx_pcs[6] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_gen3_tx_pcs[7] = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [0];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [1];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [2];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [3];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [4];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [5];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [6];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [7];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [8];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [9];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [10];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [11];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [12];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [13];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [14];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [15];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [16];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [17];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [18];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [19];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [20];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [21];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [22];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [23];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [24];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [25];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [26];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [27];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [28];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [29];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [30];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [31];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [32];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [33];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [34];
assign \w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus [35];

assign \w_hssi_gen3_tx_pcs_par_lpbk_out[0]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [0];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[1]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [1];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[2]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [2];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[3]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [3];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[4]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [4];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[5]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [5];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[6]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [6];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[7]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [7];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[8]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [8];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[9]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [9];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[10]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [10];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[11]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [11];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[12]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [12];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[13]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [13];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[14]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [14];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[15]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [15];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[16]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [16];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[17]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [17];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[18]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [18];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[19]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [19];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[20]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [20];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[21]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [21];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[22]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [22];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[23]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [23];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[24]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [24];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[25]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [25];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[26]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [26];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[27]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [27];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[28]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [28];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[29]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [29];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[30]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [30];
assign \w_hssi_gen3_tx_pcs_par_lpbk_out[31]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus [31];

assign \w_hssi_gen3_tx_pcs_tx_test_out[0]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [0];
assign \w_hssi_gen3_tx_pcs_tx_test_out[1]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [1];
assign \w_hssi_gen3_tx_pcs_tx_test_out[2]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [2];
assign \w_hssi_gen3_tx_pcs_tx_test_out[3]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [3];
assign \w_hssi_gen3_tx_pcs_tx_test_out[4]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [4];
assign \w_hssi_gen3_tx_pcs_tx_test_out[5]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [5];
assign \w_hssi_gen3_tx_pcs_tx_test_out[6]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [6];
assign \w_hssi_gen3_tx_pcs_tx_test_out[7]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [7];
assign \w_hssi_gen3_tx_pcs_tx_test_out[8]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [8];
assign \w_hssi_gen3_tx_pcs_tx_test_out[9]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [9];
assign \w_hssi_gen3_tx_pcs_tx_test_out[10]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [10];
assign \w_hssi_gen3_tx_pcs_tx_test_out[11]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [11];
assign \w_hssi_gen3_tx_pcs_tx_test_out[12]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [12];
assign \w_hssi_gen3_tx_pcs_tx_test_out[13]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [13];
assign \w_hssi_gen3_tx_pcs_tx_test_out[14]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [14];
assign \w_hssi_gen3_tx_pcs_tx_test_out[15]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [15];
assign \w_hssi_gen3_tx_pcs_tx_test_out[16]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [16];
assign \w_hssi_gen3_tx_pcs_tx_test_out[17]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [17];
assign \w_hssi_gen3_tx_pcs_tx_test_out[18]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [18];
assign \w_hssi_gen3_tx_pcs_tx_test_out[19]  = \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus [19];

assign out_avmmreaddata_hssi_krfec_tx_pcs[0] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_krfec_tx_pcs[1] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_krfec_tx_pcs[2] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_krfec_tx_pcs[3] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_krfec_tx_pcs[4] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_krfec_tx_pcs[5] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_krfec_tx_pcs[6] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_krfec_tx_pcs[7] = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_krfec_tx_pcs_tx_test_data[0]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [0];
assign \w_hssi_krfec_tx_pcs_tx_test_data[1]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [1];
assign \w_hssi_krfec_tx_pcs_tx_test_data[2]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [2];
assign \w_hssi_krfec_tx_pcs_tx_test_data[3]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [3];
assign \w_hssi_krfec_tx_pcs_tx_test_data[4]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [4];
assign \w_hssi_krfec_tx_pcs_tx_test_data[5]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [5];
assign \w_hssi_krfec_tx_pcs_tx_test_data[6]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [6];
assign \w_hssi_krfec_tx_pcs_tx_test_data[7]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [7];
assign \w_hssi_krfec_tx_pcs_tx_test_data[8]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [8];
assign \w_hssi_krfec_tx_pcs_tx_test_data[9]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [9];
assign \w_hssi_krfec_tx_pcs_tx_test_data[10]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [10];
assign \w_hssi_krfec_tx_pcs_tx_test_data[11]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [11];
assign \w_hssi_krfec_tx_pcs_tx_test_data[12]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [12];
assign \w_hssi_krfec_tx_pcs_tx_test_data[13]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [13];
assign \w_hssi_krfec_tx_pcs_tx_test_data[14]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [14];
assign \w_hssi_krfec_tx_pcs_tx_test_data[15]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [15];
assign \w_hssi_krfec_tx_pcs_tx_test_data[16]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [16];
assign \w_hssi_krfec_tx_pcs_tx_test_data[17]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [17];
assign \w_hssi_krfec_tx_pcs_tx_test_data[18]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [18];
assign \w_hssi_krfec_tx_pcs_tx_test_data[19]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus [19];

assign \w_hssi_krfec_tx_pcs_tx_data_out[0]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [0];
assign \w_hssi_krfec_tx_pcs_tx_data_out[1]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [1];
assign \w_hssi_krfec_tx_pcs_tx_data_out[2]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [2];
assign \w_hssi_krfec_tx_pcs_tx_data_out[3]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [3];
assign \w_hssi_krfec_tx_pcs_tx_data_out[4]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [4];
assign \w_hssi_krfec_tx_pcs_tx_data_out[5]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [5];
assign \w_hssi_krfec_tx_pcs_tx_data_out[6]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [6];
assign \w_hssi_krfec_tx_pcs_tx_data_out[7]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [7];
assign \w_hssi_krfec_tx_pcs_tx_data_out[8]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [8];
assign \w_hssi_krfec_tx_pcs_tx_data_out[9]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [9];
assign \w_hssi_krfec_tx_pcs_tx_data_out[10]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [10];
assign \w_hssi_krfec_tx_pcs_tx_data_out[11]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [11];
assign \w_hssi_krfec_tx_pcs_tx_data_out[12]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [12];
assign \w_hssi_krfec_tx_pcs_tx_data_out[13]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [13];
assign \w_hssi_krfec_tx_pcs_tx_data_out[14]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [14];
assign \w_hssi_krfec_tx_pcs_tx_data_out[15]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [15];
assign \w_hssi_krfec_tx_pcs_tx_data_out[16]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [16];
assign \w_hssi_krfec_tx_pcs_tx_data_out[17]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [17];
assign \w_hssi_krfec_tx_pcs_tx_data_out[18]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [18];
assign \w_hssi_krfec_tx_pcs_tx_data_out[19]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [19];
assign \w_hssi_krfec_tx_pcs_tx_data_out[20]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [20];
assign \w_hssi_krfec_tx_pcs_tx_data_out[21]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [21];
assign \w_hssi_krfec_tx_pcs_tx_data_out[22]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [22];
assign \w_hssi_krfec_tx_pcs_tx_data_out[23]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [23];
assign \w_hssi_krfec_tx_pcs_tx_data_out[24]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [24];
assign \w_hssi_krfec_tx_pcs_tx_data_out[25]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [25];
assign \w_hssi_krfec_tx_pcs_tx_data_out[26]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [26];
assign \w_hssi_krfec_tx_pcs_tx_data_out[27]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [27];
assign \w_hssi_krfec_tx_pcs_tx_data_out[28]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [28];
assign \w_hssi_krfec_tx_pcs_tx_data_out[29]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [29];
assign \w_hssi_krfec_tx_pcs_tx_data_out[30]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [30];
assign \w_hssi_krfec_tx_pcs_tx_data_out[31]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [31];
assign \w_hssi_krfec_tx_pcs_tx_data_out[32]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [32];
assign \w_hssi_krfec_tx_pcs_tx_data_out[33]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [33];
assign \w_hssi_krfec_tx_pcs_tx_data_out[34]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [34];
assign \w_hssi_krfec_tx_pcs_tx_data_out[35]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [35];
assign \w_hssi_krfec_tx_pcs_tx_data_out[36]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [36];
assign \w_hssi_krfec_tx_pcs_tx_data_out[37]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [37];
assign \w_hssi_krfec_tx_pcs_tx_data_out[38]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [38];
assign \w_hssi_krfec_tx_pcs_tx_data_out[39]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [39];
assign \w_hssi_krfec_tx_pcs_tx_data_out[40]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [40];
assign \w_hssi_krfec_tx_pcs_tx_data_out[41]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [41];
assign \w_hssi_krfec_tx_pcs_tx_data_out[42]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [42];
assign \w_hssi_krfec_tx_pcs_tx_data_out[43]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [43];
assign \w_hssi_krfec_tx_pcs_tx_data_out[44]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [44];
assign \w_hssi_krfec_tx_pcs_tx_data_out[45]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [45];
assign \w_hssi_krfec_tx_pcs_tx_data_out[46]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [46];
assign \w_hssi_krfec_tx_pcs_tx_data_out[47]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [47];
assign \w_hssi_krfec_tx_pcs_tx_data_out[48]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [48];
assign \w_hssi_krfec_tx_pcs_tx_data_out[49]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [49];
assign \w_hssi_krfec_tx_pcs_tx_data_out[50]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [50];
assign \w_hssi_krfec_tx_pcs_tx_data_out[51]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [51];
assign \w_hssi_krfec_tx_pcs_tx_data_out[52]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [52];
assign \w_hssi_krfec_tx_pcs_tx_data_out[53]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [53];
assign \w_hssi_krfec_tx_pcs_tx_data_out[54]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [54];
assign \w_hssi_krfec_tx_pcs_tx_data_out[55]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [55];
assign \w_hssi_krfec_tx_pcs_tx_data_out[56]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [56];
assign \w_hssi_krfec_tx_pcs_tx_data_out[57]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [57];
assign \w_hssi_krfec_tx_pcs_tx_data_out[58]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [58];
assign \w_hssi_krfec_tx_pcs_tx_data_out[59]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [59];
assign \w_hssi_krfec_tx_pcs_tx_data_out[60]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [60];
assign \w_hssi_krfec_tx_pcs_tx_data_out[61]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [61];
assign \w_hssi_krfec_tx_pcs_tx_data_out[62]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [62];
assign \w_hssi_krfec_tx_pcs_tx_data_out[63]  = \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus [63];

assign out_avmmreaddata_hssi_fifo_rx_pcs[0] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_fifo_rx_pcs[1] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_fifo_rx_pcs[2] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_fifo_rx_pcs[3] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_fifo_rx_pcs[4] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_fifo_rx_pcs[5] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_fifo_rx_pcs[6] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_fifo_rx_pcs[7] = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_fifo_rx_pcs_data_out2_10g[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [31];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[32]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [32];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[33]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [33];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[34]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [34];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[35]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [35];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[36]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [36];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[37]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [37];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[38]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [38];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[39]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [39];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[40]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [40];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[41]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [41];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[42]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [42];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[43]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [43];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[44]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [44];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[45]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [45];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[46]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [46];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[47]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [47];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[48]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [48];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[49]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [49];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[50]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [50];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[51]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [51];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[52]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [52];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[53]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [53];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[54]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [54];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[55]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [55];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[56]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [56];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[57]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [57];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[58]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [58];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[59]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [59];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[60]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [60];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[61]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [61];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[62]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [62];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[63]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [63];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[64]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [64];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[65]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [65];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[66]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [66];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[67]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [67];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[68]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [68];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[69]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [69];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[70]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [70];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[71]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [71];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[72]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [72];
assign \w_hssi_fifo_rx_pcs_data_out2_10g[73]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus [73];

assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus [31];

assign \w_hssi_fifo_rx_pcs_data_out_10g[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out_10g[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out_10g[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out_10g[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out_10g[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out_10g[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out_10g[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out_10g[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out_10g[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out_10g[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out_10g[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out_10g[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out_10g[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out_10g[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out_10g[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out_10g[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out_10g[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out_10g[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out_10g[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out_10g[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out_10g[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out_10g[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out_10g[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out_10g[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out_10g[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out_10g[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out_10g[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out_10g[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out_10g[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out_10g[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out_10g[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out_10g[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [31];
assign \w_hssi_fifo_rx_pcs_data_out_10g[32]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [32];
assign \w_hssi_fifo_rx_pcs_data_out_10g[33]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [33];
assign \w_hssi_fifo_rx_pcs_data_out_10g[34]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [34];
assign \w_hssi_fifo_rx_pcs_data_out_10g[35]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [35];
assign \w_hssi_fifo_rx_pcs_data_out_10g[36]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [36];
assign \w_hssi_fifo_rx_pcs_data_out_10g[37]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [37];
assign \w_hssi_fifo_rx_pcs_data_out_10g[38]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [38];
assign \w_hssi_fifo_rx_pcs_data_out_10g[39]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [39];
assign \w_hssi_fifo_rx_pcs_data_out_10g[40]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [40];
assign \w_hssi_fifo_rx_pcs_data_out_10g[41]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [41];
assign \w_hssi_fifo_rx_pcs_data_out_10g[42]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [42];
assign \w_hssi_fifo_rx_pcs_data_out_10g[43]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [43];
assign \w_hssi_fifo_rx_pcs_data_out_10g[44]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [44];
assign \w_hssi_fifo_rx_pcs_data_out_10g[45]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [45];
assign \w_hssi_fifo_rx_pcs_data_out_10g[46]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [46];
assign \w_hssi_fifo_rx_pcs_data_out_10g[47]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [47];
assign \w_hssi_fifo_rx_pcs_data_out_10g[48]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [48];
assign \w_hssi_fifo_rx_pcs_data_out_10g[49]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [49];
assign \w_hssi_fifo_rx_pcs_data_out_10g[50]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [50];
assign \w_hssi_fifo_rx_pcs_data_out_10g[51]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [51];
assign \w_hssi_fifo_rx_pcs_data_out_10g[52]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [52];
assign \w_hssi_fifo_rx_pcs_data_out_10g[53]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [53];
assign \w_hssi_fifo_rx_pcs_data_out_10g[54]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [54];
assign \w_hssi_fifo_rx_pcs_data_out_10g[55]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [55];
assign \w_hssi_fifo_rx_pcs_data_out_10g[56]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [56];
assign \w_hssi_fifo_rx_pcs_data_out_10g[57]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [57];
assign \w_hssi_fifo_rx_pcs_data_out_10g[58]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [58];
assign \w_hssi_fifo_rx_pcs_data_out_10g[59]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [59];
assign \w_hssi_fifo_rx_pcs_data_out_10g[60]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [60];
assign \w_hssi_fifo_rx_pcs_data_out_10g[61]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [61];
assign \w_hssi_fifo_rx_pcs_data_out_10g[62]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [62];
assign \w_hssi_fifo_rx_pcs_data_out_10g[63]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [63];
assign \w_hssi_fifo_rx_pcs_data_out_10g[64]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [64];
assign \w_hssi_fifo_rx_pcs_data_out_10g[65]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [65];
assign \w_hssi_fifo_rx_pcs_data_out_10g[66]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [66];
assign \w_hssi_fifo_rx_pcs_data_out_10g[67]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [67];
assign \w_hssi_fifo_rx_pcs_data_out_10g[68]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [68];
assign \w_hssi_fifo_rx_pcs_data_out_10g[69]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [69];
assign \w_hssi_fifo_rx_pcs_data_out_10g[70]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [70];
assign \w_hssi_fifo_rx_pcs_data_out_10g[71]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [71];
assign \w_hssi_fifo_rx_pcs_data_out_10g[72]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [72];
assign \w_hssi_fifo_rx_pcs_data_out_10g[73]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus [73];

assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus [31];

assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [31];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [32];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [33];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [34];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [35];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [36];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [37];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [38];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [39];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [40];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [41];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [42];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [43];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [44];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [45];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [46];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [47];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [48];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [49];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [50];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [51];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [52];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [53];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [54];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [55];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [56];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [57];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [58];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [59];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [60];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [61];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [62];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [63];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [64];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [65];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [66];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [67];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [68];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [69];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [70];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [71];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [72];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [73];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [74];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [75];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [76];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [77];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [78];
assign \w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus [79];

assign \w_hssi_fifo_rx_pcs_data_out_gen3[0]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [0];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[1]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [1];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[2]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [2];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[3]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [3];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[4]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [4];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[5]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [5];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[6]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [6];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[7]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [7];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[8]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [8];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[9]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [9];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[10]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [10];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[11]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [11];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[12]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [12];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[13]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [13];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[14]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [14];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[15]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [15];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[16]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [16];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[17]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [17];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[18]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [18];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[19]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [19];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[20]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [20];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[21]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [21];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[22]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [22];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[23]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [23];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[24]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [24];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[25]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [25];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[26]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [26];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[27]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [27];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[28]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [28];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[29]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [29];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[30]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [30];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[31]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [31];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[32]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [32];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[33]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [33];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[34]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [34];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[35]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [35];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[36]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [36];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[37]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [37];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[38]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [38];
assign \w_hssi_fifo_rx_pcs_data_out_gen3[39]  = \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus [39];

assign out_avmmreaddata_hssi_fifo_tx_pcs[0] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_fifo_tx_pcs[1] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_fifo_tx_pcs[2] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_fifo_tx_pcs[3] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_fifo_tx_pcs[4] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_fifo_tx_pcs[5] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_fifo_tx_pcs[6] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_fifo_tx_pcs[7] = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus [7];

assign \w_hssi_fifo_tx_pcs_data_out_10g[0]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [0];
assign \w_hssi_fifo_tx_pcs_data_out_10g[1]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [1];
assign \w_hssi_fifo_tx_pcs_data_out_10g[2]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [2];
assign \w_hssi_fifo_tx_pcs_data_out_10g[3]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [3];
assign \w_hssi_fifo_tx_pcs_data_out_10g[4]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [4];
assign \w_hssi_fifo_tx_pcs_data_out_10g[5]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [5];
assign \w_hssi_fifo_tx_pcs_data_out_10g[6]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [6];
assign \w_hssi_fifo_tx_pcs_data_out_10g[7]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [7];
assign \w_hssi_fifo_tx_pcs_data_out_10g[8]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [8];
assign \w_hssi_fifo_tx_pcs_data_out_10g[9]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [9];
assign \w_hssi_fifo_tx_pcs_data_out_10g[10]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [10];
assign \w_hssi_fifo_tx_pcs_data_out_10g[11]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [11];
assign \w_hssi_fifo_tx_pcs_data_out_10g[12]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [12];
assign \w_hssi_fifo_tx_pcs_data_out_10g[13]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [13];
assign \w_hssi_fifo_tx_pcs_data_out_10g[14]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [14];
assign \w_hssi_fifo_tx_pcs_data_out_10g[15]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [15];
assign \w_hssi_fifo_tx_pcs_data_out_10g[16]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [16];
assign \w_hssi_fifo_tx_pcs_data_out_10g[17]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [17];
assign \w_hssi_fifo_tx_pcs_data_out_10g[18]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [18];
assign \w_hssi_fifo_tx_pcs_data_out_10g[19]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [19];
assign \w_hssi_fifo_tx_pcs_data_out_10g[20]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [20];
assign \w_hssi_fifo_tx_pcs_data_out_10g[21]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [21];
assign \w_hssi_fifo_tx_pcs_data_out_10g[22]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [22];
assign \w_hssi_fifo_tx_pcs_data_out_10g[23]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [23];
assign \w_hssi_fifo_tx_pcs_data_out_10g[24]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [24];
assign \w_hssi_fifo_tx_pcs_data_out_10g[25]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [25];
assign \w_hssi_fifo_tx_pcs_data_out_10g[26]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [26];
assign \w_hssi_fifo_tx_pcs_data_out_10g[27]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [27];
assign \w_hssi_fifo_tx_pcs_data_out_10g[28]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [28];
assign \w_hssi_fifo_tx_pcs_data_out_10g[29]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [29];
assign \w_hssi_fifo_tx_pcs_data_out_10g[30]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [30];
assign \w_hssi_fifo_tx_pcs_data_out_10g[31]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [31];
assign \w_hssi_fifo_tx_pcs_data_out_10g[32]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [32];
assign \w_hssi_fifo_tx_pcs_data_out_10g[33]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [33];
assign \w_hssi_fifo_tx_pcs_data_out_10g[34]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [34];
assign \w_hssi_fifo_tx_pcs_data_out_10g[35]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [35];
assign \w_hssi_fifo_tx_pcs_data_out_10g[36]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [36];
assign \w_hssi_fifo_tx_pcs_data_out_10g[37]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [37];
assign \w_hssi_fifo_tx_pcs_data_out_10g[38]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [38];
assign \w_hssi_fifo_tx_pcs_data_out_10g[39]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [39];
assign \w_hssi_fifo_tx_pcs_data_out_10g[40]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [40];
assign \w_hssi_fifo_tx_pcs_data_out_10g[41]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [41];
assign \w_hssi_fifo_tx_pcs_data_out_10g[42]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [42];
assign \w_hssi_fifo_tx_pcs_data_out_10g[43]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [43];
assign \w_hssi_fifo_tx_pcs_data_out_10g[44]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [44];
assign \w_hssi_fifo_tx_pcs_data_out_10g[45]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [45];
assign \w_hssi_fifo_tx_pcs_data_out_10g[46]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [46];
assign \w_hssi_fifo_tx_pcs_data_out_10g[47]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [47];
assign \w_hssi_fifo_tx_pcs_data_out_10g[48]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [48];
assign \w_hssi_fifo_tx_pcs_data_out_10g[49]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [49];
assign \w_hssi_fifo_tx_pcs_data_out_10g[50]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [50];
assign \w_hssi_fifo_tx_pcs_data_out_10g[51]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [51];
assign \w_hssi_fifo_tx_pcs_data_out_10g[52]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [52];
assign \w_hssi_fifo_tx_pcs_data_out_10g[53]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [53];
assign \w_hssi_fifo_tx_pcs_data_out_10g[54]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [54];
assign \w_hssi_fifo_tx_pcs_data_out_10g[55]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [55];
assign \w_hssi_fifo_tx_pcs_data_out_10g[56]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [56];
assign \w_hssi_fifo_tx_pcs_data_out_10g[57]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [57];
assign \w_hssi_fifo_tx_pcs_data_out_10g[58]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [58];
assign \w_hssi_fifo_tx_pcs_data_out_10g[59]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [59];
assign \w_hssi_fifo_tx_pcs_data_out_10g[60]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [60];
assign \w_hssi_fifo_tx_pcs_data_out_10g[61]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [61];
assign \w_hssi_fifo_tx_pcs_data_out_10g[62]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [62];
assign \w_hssi_fifo_tx_pcs_data_out_10g[63]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [63];
assign \w_hssi_fifo_tx_pcs_data_out_10g[64]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [64];
assign \w_hssi_fifo_tx_pcs_data_out_10g[65]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [65];
assign \w_hssi_fifo_tx_pcs_data_out_10g[66]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [66];
assign \w_hssi_fifo_tx_pcs_data_out_10g[67]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [67];
assign \w_hssi_fifo_tx_pcs_data_out_10g[68]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [68];
assign \w_hssi_fifo_tx_pcs_data_out_10g[69]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [69];
assign \w_hssi_fifo_tx_pcs_data_out_10g[70]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [70];
assign \w_hssi_fifo_tx_pcs_data_out_10g[71]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [71];
assign \w_hssi_fifo_tx_pcs_data_out_10g[72]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus [72];

assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [0];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [1];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [2];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [3];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [4];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [5];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [6];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [7];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [8];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [9];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [10];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [11];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [12];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [13];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [14];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [15];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [16];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [17];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [18];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [19];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [20];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [21];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [22];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [23];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [24];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [25];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [26];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [27];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [28];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [29];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [30];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [31];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [32];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [33];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [34];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [35];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [36];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [37];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [38];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [39];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [40];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [41];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [42];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [43];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [44];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [45];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [46];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [47];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [48];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [49];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [50];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [51];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [52];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [53];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [54];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [55];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [56];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [57];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [58];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [59];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [60];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [61];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [62];
assign \w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63]  = \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus [63];

assign out_avmmreaddata_hssi_common_pcs_pma_interface[0] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[1] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[2] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[3] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[4] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[5] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[6] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_common_pcs_pma_interface[7] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus [7];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [2];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [3];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [4];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [5];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [7];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus [8];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [1];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [2];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [3];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [4];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [5];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [6];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [7];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus [8];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PCIE_SW_DONE_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PCIE_SW_DONE_bus [1];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus [1];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus [2];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus [3];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus [4];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [1];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [2];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [3];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [4];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [5];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [6];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [7];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [8];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [9];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [10];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [11];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [12];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [13];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [14];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [15];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [16];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [17];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [18];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus [19];

assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [0];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [1];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [2];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [3];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [4];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [5];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [6];
assign \w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7]  = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus [7];

assign out_pma_current_coeff[0] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [0];
assign out_pma_current_coeff[1] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [1];
assign out_pma_current_coeff[2] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [2];
assign out_pma_current_coeff[3] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [3];
assign out_pma_current_coeff[4] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [4];
assign out_pma_current_coeff[5] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [5];
assign out_pma_current_coeff[6] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [6];
assign out_pma_current_coeff[7] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [7];
assign out_pma_current_coeff[8] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [8];
assign out_pma_current_coeff[9] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [9];
assign out_pma_current_coeff[10] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [10];
assign out_pma_current_coeff[11] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [11];
assign out_pma_current_coeff[12] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [12];
assign out_pma_current_coeff[13] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [13];
assign out_pma_current_coeff[14] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [14];
assign out_pma_current_coeff[15] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [15];
assign out_pma_current_coeff[16] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [16];
assign out_pma_current_coeff[17] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus [17];

assign out_pma_pcie_switch[0] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_PCIE_SWITCH_bus [0];
assign out_pma_pcie_switch[1] = \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_PCIE_SWITCH_bus [1];

assign out_avmmreaddata_hssi_tx_pcs_pma_interface[0] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [0];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[1] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [1];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[2] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [2];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[3] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [3];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[4] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [4];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[5] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [5];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[6] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [6];
assign out_avmmreaddata_hssi_tx_pcs_pma_interface[7] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus [7];

assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT0  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [0];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT1  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [1];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT2  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [2];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT3  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [3];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT4  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [4];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT5  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [5];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT6  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [6];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT7  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [7];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT8  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [8];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT9  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [9];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT10  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [10];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT11  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [11];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT12  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [12];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT13  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [13];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT14  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [14];
assign \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface~O_AVMM_USER_DATAOUT15  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus [15];

assign \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus [0];
assign \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus [1];
assign \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus [2];
assign \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus [3];
assign \w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus [4];

assign out_pma_tx_pma_data[0] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [0];
assign out_pma_tx_pma_data[1] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [1];
assign out_pma_tx_pma_data[2] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [2];
assign out_pma_tx_pma_data[3] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [3];
assign out_pma_tx_pma_data[4] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [4];
assign out_pma_tx_pma_data[5] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [5];
assign out_pma_tx_pma_data[6] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [6];
assign out_pma_tx_pma_data[7] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [7];
assign out_pma_tx_pma_data[8] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [8];
assign out_pma_tx_pma_data[9] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [9];
assign out_pma_tx_pma_data[10] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [10];
assign out_pma_tx_pma_data[11] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [11];
assign out_pma_tx_pma_data[12] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [12];
assign out_pma_tx_pma_data[13] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [13];
assign out_pma_tx_pma_data[14] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [14];
assign out_pma_tx_pma_data[15] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [15];
assign out_pma_tx_pma_data[16] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [16];
assign out_pma_tx_pma_data[17] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [17];
assign out_pma_tx_pma_data[18] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [18];
assign out_pma_tx_pma_data[19] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [19];
assign out_pma_tx_pma_data[20] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [20];
assign out_pma_tx_pma_data[21] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [21];
assign out_pma_tx_pma_data[22] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [22];
assign out_pma_tx_pma_data[23] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [23];
assign out_pma_tx_pma_data[24] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [24];
assign out_pma_tx_pma_data[25] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [25];
assign out_pma_tx_pma_data[26] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [26];
assign out_pma_tx_pma_data[27] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [27];
assign out_pma_tx_pma_data[28] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [28];
assign out_pma_tx_pma_data[29] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [29];
assign out_pma_tx_pma_data[30] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [30];
assign out_pma_tx_pma_data[31] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [31];
assign out_pma_tx_pma_data[32] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [32];
assign out_pma_tx_pma_data[33] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [33];
assign out_pma_tx_pma_data[34] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [34];
assign out_pma_tx_pma_data[35] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [35];
assign out_pma_tx_pma_data[36] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [36];
assign out_pma_tx_pma_data[37] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [37];
assign out_pma_tx_pma_data[38] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [38];
assign out_pma_tx_pma_data[39] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [39];
assign out_pma_tx_pma_data[40] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [40];
assign out_pma_tx_pma_data[41] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [41];
assign out_pma_tx_pma_data[42] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [42];
assign out_pma_tx_pma_data[43] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [43];
assign out_pma_tx_pma_data[44] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [44];
assign out_pma_tx_pma_data[45] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [45];
assign out_pma_tx_pma_data[46] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [46];
assign out_pma_tx_pma_data[47] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [47];
assign out_pma_tx_pma_data[48] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [48];
assign out_pma_tx_pma_data[49] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [49];
assign out_pma_tx_pma_data[50] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [50];
assign out_pma_tx_pma_data[51] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [51];
assign out_pma_tx_pma_data[52] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [52];
assign out_pma_tx_pma_data[53] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [53];
assign out_pma_tx_pma_data[54] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [54];
assign out_pma_tx_pma_data[55] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [55];
assign out_pma_tx_pma_data[56] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [56];
assign out_pma_tx_pma_data[57] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [57];
assign out_pma_tx_pma_data[58] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [58];
assign out_pma_tx_pma_data[59] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [59];
assign out_pma_tx_pma_data[60] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [60];
assign out_pma_tx_pma_data[61] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [61];
assign out_pma_tx_pma_data[62] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [62];
assign out_pma_tx_pma_data[63] = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus [63];

assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [0];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [1];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [2];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [3];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [4];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [5];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [6];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [7];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [8];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [9];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [10];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [11];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [12];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [13];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [14];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [15];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [16];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [17];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [18];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [19];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [20];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [21];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [22];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [23];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [24];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [25];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [26];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [27];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [28];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [29];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [30];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [31];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [32];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [33];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [34];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [35];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [36];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [37];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [38];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [39];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [40];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [41];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [42];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [43];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [44];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [45];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [46];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [47];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [48];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [49];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [50];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [51];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [52];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [53];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [54];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [55];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [56];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [57];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [58];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [59];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [60];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [61];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [62];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus [63];

assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [0];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [1];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [2];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [3];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [4];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [5];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [6];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [7];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [8];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [9];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [10];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [11];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [12];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [13];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [14];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [15];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [16];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [17];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [18];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [19];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [20];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [21];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [22];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [23];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [24];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [25];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [26];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [27];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [28];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [29];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [30];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [31];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [32];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [33];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [34];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [35];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [36];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [37];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [38];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [39];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [40];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [41];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [42];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [43];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [44];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [45];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [46];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [47];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [48];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [49];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [50];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [51];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [52];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [53];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [54];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [55];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [56];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [57];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [58];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [59];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [60];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [61];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [62];
assign \w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus [63];

assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [0];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [1];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [2];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [3];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [4];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [5];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [6];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [7];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [8];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [9];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [10];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [11];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [12];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [13];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [14];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [15];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [16];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [17];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [18];
assign \w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus [19];

assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [0];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [1];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [2];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [3];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [4];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [5];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [6];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [7];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [8];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [9];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [10];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [11];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [12];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [13];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [14];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [15];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [16];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [17];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [18];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus [19];

assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [0];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [1];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [2];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [3];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [4];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [5];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [6];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [7];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [8];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [9];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [10];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [11];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [12];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [13];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [14];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [15];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [16];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [17];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [18];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus [19];

assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [0];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [1];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [2];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [3];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [4];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [5];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [6];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [7];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [8];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [9];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [10];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [11];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [12];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [13];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [14];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [15];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [16];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [17];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [18];
assign \w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19]  = \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus [19];

twentynm_hssi_rx_pld_pcs_interface \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pldif_10g_rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
	.int_pldif_10g_rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
	.int_pldif_10g_rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
	.int_pldif_10g_rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
	.int_pldif_10g_rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
	.int_pldif_10g_rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
	.int_pldif_10g_rx_empty(w_hssi_10g_rx_pcs_rx_empty),
	.int_pldif_10g_rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
	.int_pldif_10g_rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
	.int_pldif_10g_rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
	.int_pldif_10g_rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
	.int_pldif_10g_rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
	.int_pldif_10g_rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
	.int_pldif_10g_rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
	.int_pldif_10g_rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
	.int_pldif_8g_empty_rmf(w_hssi_8g_rx_pcs_rm_fifo_empty),
	.int_pldif_8g_empty_rx(w_hssi_8g_rx_pcs_pc_fifo_empty),
	.int_pldif_8g_full_rmf(w_hssi_8g_rx_pcs_rm_fifo_full),
	.int_pldif_8g_full_rx(w_hssi_8g_rx_pcs_pcfifofull),
	.int_pldif_8g_phystatus(w_hssi_8g_rx_pcs_phystatus),
	.int_pldif_8g_rx_clk(w_hssi_8g_rx_pcs_clock_to_pld),
	.int_pldif_8g_rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
	.int_pldif_8g_rx_rstn_sync2wrfifo(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
	.int_pldif_8g_rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
	.int_pldif_8g_rxvalid(w_hssi_8g_rx_pcs_rxvalid),
	.int_pldif_8g_signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
	.int_pldif_krfec_rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
	.int_pldif_krfec_rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
	.int_pldif_pmaif_clkdiv_rx(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
	.int_pldif_pmaif_clkdiv_rx_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
	.int_pldif_pmaif_rx_prbs_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
	.int_pldif_pmaif_rx_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
	.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
	.int_pldif_pmaif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
	.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
	.pld_10g_krfec_rx_clr_errblk_cnt(gnd),
	.pld_10g_krfec_rx_pld_rst_n(!in_pld_10g_krfec_rx_pld_rst_n),
	.pld_10g_rx_align_clr(gnd),
	.pld_10g_rx_clr_ber_count(gnd),
	.pld_10g_rx_rd_en(gnd),
	.pld_8g_a1a2_size(gnd),
	.pld_8g_bitloc_rev_en(gnd),
	.pld_8g_byte_rev_en(gnd),
	.pld_8g_encdt(in_pld_8g_encdt),
	.pld_8g_g3_rx_pld_rst_n(!in_pld_10g_krfec_rx_pld_rst_n),
	.pld_8g_rdenable_rx(gnd),
	.pld_8g_rxpolarity(gnd),
	.pld_8g_wrdisable_rx(gnd),
	.pld_bitslip(gnd),
	.pld_partial_reconfig(vcc),
	.pld_pma_rxpma_rstb(!in_pld_pma_rxpma_rstb),
	.pld_pmaif_rx_pld_rst_n(!in_pld_10g_krfec_rx_pld_rst_n),
	.pld_pmaif_rxclkslip(gnd),
	.pld_polinv_rx(gnd),
	.pld_rx_clk(in_pld_rx_clk),
	.pld_rx_prbs_err_clr(gnd),
	.pld_syncsm_en(vcc),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.int_pldif_10g_rx_control({\w_hssi_10g_rx_pcs_rx_control[19] ,\w_hssi_10g_rx_pcs_rx_control[18] ,\w_hssi_10g_rx_pcs_rx_control[17] ,\w_hssi_10g_rx_pcs_rx_control[16] ,\w_hssi_10g_rx_pcs_rx_control[15] ,\w_hssi_10g_rx_pcs_rx_control[14] ,\w_hssi_10g_rx_pcs_rx_control[13] ,
\w_hssi_10g_rx_pcs_rx_control[12] ,\w_hssi_10g_rx_pcs_rx_control[11] ,\w_hssi_10g_rx_pcs_rx_control[10] ,\w_hssi_10g_rx_pcs_rx_control[9] ,\w_hssi_10g_rx_pcs_rx_control[8] ,\w_hssi_10g_rx_pcs_rx_control[7] ,\w_hssi_10g_rx_pcs_rx_control[6] ,
\w_hssi_10g_rx_pcs_rx_control[5] ,\w_hssi_10g_rx_pcs_rx_control[4] ,\w_hssi_10g_rx_pcs_rx_control[3] ,\w_hssi_10g_rx_pcs_rx_control[2] ,\w_hssi_10g_rx_pcs_rx_control[1] ,\w_hssi_10g_rx_pcs_rx_control[0] }),
	.int_pldif_10g_rx_data({\w_hssi_10g_rx_pcs_rx_data[127] ,\w_hssi_10g_rx_pcs_rx_data[126] ,\w_hssi_10g_rx_pcs_rx_data[125] ,\w_hssi_10g_rx_pcs_rx_data[124] ,\w_hssi_10g_rx_pcs_rx_data[123] ,\w_hssi_10g_rx_pcs_rx_data[122] ,\w_hssi_10g_rx_pcs_rx_data[121] ,\w_hssi_10g_rx_pcs_rx_data[120] ,
\w_hssi_10g_rx_pcs_rx_data[119] ,\w_hssi_10g_rx_pcs_rx_data[118] ,\w_hssi_10g_rx_pcs_rx_data[117] ,\w_hssi_10g_rx_pcs_rx_data[116] ,\w_hssi_10g_rx_pcs_rx_data[115] ,\w_hssi_10g_rx_pcs_rx_data[114] ,\w_hssi_10g_rx_pcs_rx_data[113] ,\w_hssi_10g_rx_pcs_rx_data[112] ,
\w_hssi_10g_rx_pcs_rx_data[111] ,\w_hssi_10g_rx_pcs_rx_data[110] ,\w_hssi_10g_rx_pcs_rx_data[109] ,\w_hssi_10g_rx_pcs_rx_data[108] ,\w_hssi_10g_rx_pcs_rx_data[107] ,\w_hssi_10g_rx_pcs_rx_data[106] ,\w_hssi_10g_rx_pcs_rx_data[105] ,\w_hssi_10g_rx_pcs_rx_data[104] ,
\w_hssi_10g_rx_pcs_rx_data[103] ,\w_hssi_10g_rx_pcs_rx_data[102] ,\w_hssi_10g_rx_pcs_rx_data[101] ,\w_hssi_10g_rx_pcs_rx_data[100] ,\w_hssi_10g_rx_pcs_rx_data[99] ,\w_hssi_10g_rx_pcs_rx_data[98] ,\w_hssi_10g_rx_pcs_rx_data[97] ,\w_hssi_10g_rx_pcs_rx_data[96] ,
\w_hssi_10g_rx_pcs_rx_data[95] ,\w_hssi_10g_rx_pcs_rx_data[94] ,\w_hssi_10g_rx_pcs_rx_data[93] ,\w_hssi_10g_rx_pcs_rx_data[92] ,\w_hssi_10g_rx_pcs_rx_data[91] ,\w_hssi_10g_rx_pcs_rx_data[90] ,\w_hssi_10g_rx_pcs_rx_data[89] ,\w_hssi_10g_rx_pcs_rx_data[88] ,
\w_hssi_10g_rx_pcs_rx_data[87] ,\w_hssi_10g_rx_pcs_rx_data[86] ,\w_hssi_10g_rx_pcs_rx_data[85] ,\w_hssi_10g_rx_pcs_rx_data[84] ,\w_hssi_10g_rx_pcs_rx_data[83] ,\w_hssi_10g_rx_pcs_rx_data[82] ,\w_hssi_10g_rx_pcs_rx_data[81] ,\w_hssi_10g_rx_pcs_rx_data[80] ,
\w_hssi_10g_rx_pcs_rx_data[79] ,\w_hssi_10g_rx_pcs_rx_data[78] ,\w_hssi_10g_rx_pcs_rx_data[77] ,\w_hssi_10g_rx_pcs_rx_data[76] ,\w_hssi_10g_rx_pcs_rx_data[75] ,\w_hssi_10g_rx_pcs_rx_data[74] ,\w_hssi_10g_rx_pcs_rx_data[73] ,\w_hssi_10g_rx_pcs_rx_data[72] ,
\w_hssi_10g_rx_pcs_rx_data[71] ,\w_hssi_10g_rx_pcs_rx_data[70] ,\w_hssi_10g_rx_pcs_rx_data[69] ,\w_hssi_10g_rx_pcs_rx_data[68] ,\w_hssi_10g_rx_pcs_rx_data[67] ,\w_hssi_10g_rx_pcs_rx_data[66] ,\w_hssi_10g_rx_pcs_rx_data[65] ,\w_hssi_10g_rx_pcs_rx_data[64] ,
\w_hssi_10g_rx_pcs_rx_data[63] ,\w_hssi_10g_rx_pcs_rx_data[62] ,\w_hssi_10g_rx_pcs_rx_data[61] ,\w_hssi_10g_rx_pcs_rx_data[60] ,\w_hssi_10g_rx_pcs_rx_data[59] ,\w_hssi_10g_rx_pcs_rx_data[58] ,\w_hssi_10g_rx_pcs_rx_data[57] ,\w_hssi_10g_rx_pcs_rx_data[56] ,
\w_hssi_10g_rx_pcs_rx_data[55] ,\w_hssi_10g_rx_pcs_rx_data[54] ,\w_hssi_10g_rx_pcs_rx_data[53] ,\w_hssi_10g_rx_pcs_rx_data[52] ,\w_hssi_10g_rx_pcs_rx_data[51] ,\w_hssi_10g_rx_pcs_rx_data[50] ,\w_hssi_10g_rx_pcs_rx_data[49] ,\w_hssi_10g_rx_pcs_rx_data[48] ,
\w_hssi_10g_rx_pcs_rx_data[47] ,\w_hssi_10g_rx_pcs_rx_data[46] ,\w_hssi_10g_rx_pcs_rx_data[45] ,\w_hssi_10g_rx_pcs_rx_data[44] ,\w_hssi_10g_rx_pcs_rx_data[43] ,\w_hssi_10g_rx_pcs_rx_data[42] ,\w_hssi_10g_rx_pcs_rx_data[41] ,\w_hssi_10g_rx_pcs_rx_data[40] ,
\w_hssi_10g_rx_pcs_rx_data[39] ,\w_hssi_10g_rx_pcs_rx_data[38] ,\w_hssi_10g_rx_pcs_rx_data[37] ,\w_hssi_10g_rx_pcs_rx_data[36] ,\w_hssi_10g_rx_pcs_rx_data[35] ,\w_hssi_10g_rx_pcs_rx_data[34] ,\w_hssi_10g_rx_pcs_rx_data[33] ,\w_hssi_10g_rx_pcs_rx_data[32] ,
\w_hssi_10g_rx_pcs_rx_data[31] ,\w_hssi_10g_rx_pcs_rx_data[30] ,\w_hssi_10g_rx_pcs_rx_data[29] ,\w_hssi_10g_rx_pcs_rx_data[28] ,\w_hssi_10g_rx_pcs_rx_data[27] ,\w_hssi_10g_rx_pcs_rx_data[26] ,\w_hssi_10g_rx_pcs_rx_data[25] ,\w_hssi_10g_rx_pcs_rx_data[24] ,
\w_hssi_10g_rx_pcs_rx_data[23] ,\w_hssi_10g_rx_pcs_rx_data[22] ,\w_hssi_10g_rx_pcs_rx_data[21] ,\w_hssi_10g_rx_pcs_rx_data[20] ,\w_hssi_10g_rx_pcs_rx_data[19] ,\w_hssi_10g_rx_pcs_rx_data[18] ,\w_hssi_10g_rx_pcs_rx_data[17] ,\w_hssi_10g_rx_pcs_rx_data[16] ,
\w_hssi_10g_rx_pcs_rx_data[15] ,\w_hssi_10g_rx_pcs_rx_data[14] ,\w_hssi_10g_rx_pcs_rx_data[13] ,\w_hssi_10g_rx_pcs_rx_data[12] ,\w_hssi_10g_rx_pcs_rx_data[11] ,\w_hssi_10g_rx_pcs_rx_data[10] ,\w_hssi_10g_rx_pcs_rx_data[9] ,\w_hssi_10g_rx_pcs_rx_data[8] ,
\w_hssi_10g_rx_pcs_rx_data[7] ,\w_hssi_10g_rx_pcs_rx_data[6] ,\w_hssi_10g_rx_pcs_rx_data[5] ,\w_hssi_10g_rx_pcs_rx_data[4] ,\w_hssi_10g_rx_pcs_rx_data[3] ,\w_hssi_10g_rx_pcs_rx_data[2] ,\w_hssi_10g_rx_pcs_rx_data[1] ,\w_hssi_10g_rx_pcs_rx_data[0] }),
	.int_pldif_10g_rx_diag_status({\w_hssi_10g_rx_pcs_rx_diag_status[1] ,\w_hssi_10g_rx_pcs_rx_diag_status[0] }),
	.int_pldif_10g_rx_fifo_num({\w_hssi_10g_rx_pcs_rx_fifo_num[4] ,\w_hssi_10g_rx_pcs_rx_fifo_num[3] ,\w_hssi_10g_rx_pcs_rx_fifo_num[2] ,\w_hssi_10g_rx_pcs_rx_fifo_num[1] ,\w_hssi_10g_rx_pcs_rx_fifo_num[0] }),
	.int_pldif_8g_a1a2_k1k2_flag({\w_hssi_8g_rx_pcs_a1a2k1k2flag[3] ,\w_hssi_8g_rx_pcs_a1a2k1k2flag[2] ,\w_hssi_8g_rx_pcs_a1a2k1k2flag[1] ,\w_hssi_8g_rx_pcs_a1a2k1k2flag[0] }),
	.int_pldif_8g_rx_blk_start({\w_hssi_8g_rx_pcs_rx_blk_start[3] ,\w_hssi_8g_rx_pcs_rx_blk_start[2] ,\w_hssi_8g_rx_pcs_rx_blk_start[1] ,\w_hssi_8g_rx_pcs_rx_blk_start[0] }),
	.int_pldif_8g_rx_data_valid({\w_hssi_8g_rx_pcs_rx_data_valid[3] ,\w_hssi_8g_rx_pcs_rx_data_valid[2] ,\w_hssi_8g_rx_pcs_rx_data_valid[1] ,\w_hssi_8g_rx_pcs_rx_data_valid[0] }),
	.int_pldif_8g_rx_sync_hdr({\w_hssi_8g_rx_pcs_rx_sync_hdr[1] ,\w_hssi_8g_rx_pcs_rx_sync_hdr[0] }),
	.int_pldif_8g_rxd({\w_hssi_8g_rx_pcs_dataout[63] ,\w_hssi_8g_rx_pcs_dataout[62] ,\w_hssi_8g_rx_pcs_dataout[61] ,\w_hssi_8g_rx_pcs_dataout[60] ,\w_hssi_8g_rx_pcs_dataout[59] ,\w_hssi_8g_rx_pcs_dataout[58] ,\w_hssi_8g_rx_pcs_dataout[57] ,\w_hssi_8g_rx_pcs_dataout[56] ,
\w_hssi_8g_rx_pcs_dataout[55] ,\w_hssi_8g_rx_pcs_dataout[54] ,\w_hssi_8g_rx_pcs_dataout[53] ,\w_hssi_8g_rx_pcs_dataout[52] ,\w_hssi_8g_rx_pcs_dataout[51] ,\w_hssi_8g_rx_pcs_dataout[50] ,\w_hssi_8g_rx_pcs_dataout[49] ,\w_hssi_8g_rx_pcs_dataout[48] ,
\w_hssi_8g_rx_pcs_dataout[47] ,\w_hssi_8g_rx_pcs_dataout[46] ,\w_hssi_8g_rx_pcs_dataout[45] ,\w_hssi_8g_rx_pcs_dataout[44] ,\w_hssi_8g_rx_pcs_dataout[43] ,\w_hssi_8g_rx_pcs_dataout[42] ,\w_hssi_8g_rx_pcs_dataout[41] ,\w_hssi_8g_rx_pcs_dataout[40] ,
\w_hssi_8g_rx_pcs_dataout[39] ,\w_hssi_8g_rx_pcs_dataout[38] ,\w_hssi_8g_rx_pcs_dataout[37] ,\w_hssi_8g_rx_pcs_dataout[36] ,\w_hssi_8g_rx_pcs_dataout[35] ,\w_hssi_8g_rx_pcs_dataout[34] ,\w_hssi_8g_rx_pcs_dataout[33] ,\w_hssi_8g_rx_pcs_dataout[32] ,
\w_hssi_8g_rx_pcs_dataout[31] ,\w_hssi_8g_rx_pcs_dataout[30] ,\w_hssi_8g_rx_pcs_dataout[29] ,\w_hssi_8g_rx_pcs_dataout[28] ,\w_hssi_8g_rx_pcs_dataout[27] ,\w_hssi_8g_rx_pcs_dataout[26] ,\w_hssi_8g_rx_pcs_dataout[25] ,\w_hssi_8g_rx_pcs_dataout[24] ,
\w_hssi_8g_rx_pcs_dataout[23] ,\w_hssi_8g_rx_pcs_dataout[22] ,\w_hssi_8g_rx_pcs_dataout[21] ,\w_hssi_8g_rx_pcs_dataout[20] ,\w_hssi_8g_rx_pcs_dataout[19] ,\w_hssi_8g_rx_pcs_dataout[18] ,\w_hssi_8g_rx_pcs_dataout[17] ,\w_hssi_8g_rx_pcs_dataout[16] ,
\w_hssi_8g_rx_pcs_dataout[15] ,\w_hssi_8g_rx_pcs_dataout[14] ,\w_hssi_8g_rx_pcs_dataout[13] ,\w_hssi_8g_rx_pcs_dataout[12] ,\w_hssi_8g_rx_pcs_dataout[11] ,\w_hssi_8g_rx_pcs_dataout[10] ,\w_hssi_8g_rx_pcs_dataout[9] ,\w_hssi_8g_rx_pcs_dataout[8] ,
\w_hssi_8g_rx_pcs_dataout[7] ,\w_hssi_8g_rx_pcs_dataout[6] ,\w_hssi_8g_rx_pcs_dataout[5] ,\w_hssi_8g_rx_pcs_dataout[4] ,\w_hssi_8g_rx_pcs_dataout[3] ,\w_hssi_8g_rx_pcs_dataout[2] ,\w_hssi_8g_rx_pcs_dataout[1] ,\w_hssi_8g_rx_pcs_dataout[0] }),
	.int_pldif_8g_rxstatus({\w_hssi_8g_rx_pcs_rxstatus[2] ,\w_hssi_8g_rx_pcs_rxstatus[1] ,\w_hssi_8g_rx_pcs_rxstatus[0] }),
	.int_pldif_8g_wa_boundary({\w_hssi_8g_rx_pcs_word_align_boundary[4] ,\w_hssi_8g_rx_pcs_word_align_boundary[3] ,\w_hssi_8g_rx_pcs_word_align_boundary[2] ,\w_hssi_8g_rx_pcs_word_align_boundary[1] ,\w_hssi_8g_rx_pcs_word_align_boundary[0] }),
	.int_pldif_krfec_rx_data_status({\w_hssi_krfec_rx_pcs_rx_data_status[1] ,\w_hssi_krfec_rx_pcs_rx_data_status[0] }),
	.int_pldif_pmaif_rx_data({\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[63] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[62] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[61] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[60] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[59] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[58] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[57] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[56] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[55] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[54] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[53] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[52] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[51] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[50] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[49] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[48] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[47] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[46] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[45] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[44] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[43] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[42] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[41] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[40] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[39] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[38] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[37] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[36] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[35] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[34] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[33] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[32] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[31] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[30] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[29] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[28] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[27] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[26] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[25] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[24] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[23] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[22] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[21] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[20] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[19] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[18] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[17] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[16] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[15] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[14] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[13] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[12] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[11] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[10] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[9] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[8] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[7] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[6] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[5] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[4] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[3] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[2] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[1] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_data[0] }),
	.blockselect(out_blockselect_hssi_rx_pld_pcs_interface),
	.int_pldif_10g_rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
	.int_pldif_10g_rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
	.int_pldif_10g_rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
	.int_pldif_10g_rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
	.int_pldif_10g_rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
	.int_pldif_10g_rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
	.int_pldif_10g_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
	.int_pldif_10g_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
	.int_pldif_10g_rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
	.int_pldif_8g_a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
	.int_pldif_8g_bitloc_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
	.int_pldif_8g_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
	.int_pldif_8g_byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
	.int_pldif_8g_encdt(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
	.int_pldif_8g_pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
	.int_pldif_8g_rdenable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
	.int_pldif_8g_rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
	.int_pldif_8g_rxurstpcs_n(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
	.int_pldif_8g_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
	.int_pldif_8g_wrdisable_rx(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
	.int_pldif_g3_syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
	.int_pldif_krfec_rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
	.int_pldif_pmaif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
	.int_pldif_pmaif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
	.int_pldif_pmaif_rx_pld_clk(),
	.int_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
	.int_pldif_pmaif_rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
	.int_pldif_pmaif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
	.pld_10g_krfec_rx_blk_lock(),
	.pld_10g_krfec_rx_frame(),
	.pld_10g_rx_align_val(),
	.pld_10g_rx_crc32_err(),
	.pld_10g_rx_data_valid(),
	.pld_10g_rx_empty(),
	.pld_10g_rx_fifo_del(),
	.pld_10g_rx_fifo_insert(),
	.pld_10g_rx_frame_lock(),
	.pld_10g_rx_hi_ber(),
	.pld_10g_rx_oflw_err(),
	.pld_10g_rx_pempty(),
	.pld_10g_rx_pfull(),
	.pld_8g_empty_rmf(),
	.pld_8g_empty_rx(),
	.pld_8g_full_rmf(),
	.pld_8g_full_rx(),
	.pld_8g_rxelecidle(),
	.pld_8g_signal_detect_out(),
	.pld_8g_wa_boundary_txclk_fastreg(),
	.pld_8g_wa_boundary_txclk_reg(),
	.pld_bitslip_10g_txclk_reg(),
	.pld_bitslip_8g_txclk_reg(),
	.pld_bitslip_rxclk_parallel_loopback_reg(),
	.pld_bitslip_rxclk_reg(),
	.pld_pcs_rx_clk_out(out_pld_pcs_rx_clk_out),
	.pld_pcs_rx_clk_out_pcsdirect_wire(),
	.pld_pma_clkdiv_rx_user(),
	.pld_pma_rx_clk_out(),
	.pld_pma_rx_clk_out_10g_or_pcsdirect_wire(),
	.pld_pma_rx_clk_out_8g_wire(),
	.pld_pma_signal_ok(),
	.pld_pmaif_rx_pld_rst_n_reg(),
	.pld_pmaif_tx_pld_rst_n_txclk_reg(),
	.pld_polinv_rx_reg(),
	.pld_rx_clk_fifo(),
	.pld_rx_control_fifo(),
	.pld_rx_control_pcsdirect_reg(),
	.pld_rx_data_fifo(),
	.pld_rx_data_pcsdirect_reg(),
	.pld_rx_prbs_done(),
	.pld_rx_prbs_done_reg(),
	.pld_rx_prbs_done_txclk_reg(),
	.pld_rx_prbs_err(),
	.pld_rx_prbs_err_clr_pcsdirect_txclk_reg(),
	.pld_rx_prbs_err_clr_reg(),
	.pld_rx_prbs_err_disprbs_reg(),
	.pld_rx_prbs_err_pcsdirect_txclk_reg(),
	.pld_rx_prbs_err_reg(),
	.pma_rx_pma_clk_reg(),
	.avmmreaddata(\gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_AVMMREADDATA_bus ),
	.hip_rx_ctrl(),
	.hip_rx_data(),
	.int_pldif_10g_rx_control_fb(\gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_CONTROL_FB_bus ),
	.int_pldif_10g_rx_data_fb(\gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_INT_PLDIF_10G_RX_DATA_FB_bus ),
	.pld_10g_krfec_rx_diag_data_status(),
	.pld_10g_rx_fifo_num(),
	.pld_8g_a1a2_k1k2_flag(),
	.pld_8g_wa_boundary(\gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_8G_WA_BOUNDARY_bus ),
	.pld_rx_control(),
	.pld_rx_data(\gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface_PLD_RX_DATA_bus ));
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_advanced_user_mode_rx = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_ctrl_plane_bonding_rx = "individual_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_fifo_mode_rx = "fifo_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_low_latency_en_rx = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_pma_dw_rx = "pma_64b_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_prot_mode_rx = "disabled_prot_mode_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_shared_fifo_width_rx = "single_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_10g_test_bus_mode = "rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_ctrl_plane_bonding_rx = "individual_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_fifo_mode_rx = "reg_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_hip_mode = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_pma_dw_rx = "pma_10b_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_prot_mode_rx = "cpri_rx_tx_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_8g_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_clklow_clk_hz = 30'b000111011100110101100101000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_ctrl_plane_bonding_rx = "individual_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_fref_clk_hz = 30'b000111011100110101100101000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_frequency_rules_en = "enable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_func_mode = "enable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_hclk_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_hip_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_hrdrstctl_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_low_latency_en_rx = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_operating_voltage = "standard";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pcs_ac_pwr_rules_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pcs_pair_ac_pwr_uw_per_mhz = 20'b00000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pcs_rx_ac_pwr_uw_per_mhz = 20'b00000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pcs_rx_pwr_scaling_clk = "pma_rx_clk";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pld_fifo_mode_rx = "reg_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pld_rx_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pma_dw_rx = "pma_10b_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_pma_rx_clk_hz = 30'b000111011100110101100101000000;
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_prot_mode_rx = "cpri_8b10b_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_shared_fifo_width_rx = "single_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_speed_grade = "e2";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_chnl_transparent_pcs_rx = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_fifo_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_fifo_prot_mode_rx = "non_teng_mode_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_fifo_shared_fifo_width_rx = "single_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_fifo_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_g3_prot_mode = "disabled_prot_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_g3_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_low_latency_en_rx = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_prot_mode_rx = "disabled_prot_mode_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_krfec_test_bus_mode = "tx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pldif_hrdrstctl_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pldif_prot_mode_rx = "eightg_and_g3_reg_mode_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pldif_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_pma_dw_rx = "pma_10b_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_prot_mode_rx = "eightg_only_pld_mode_rx";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_sim_mode = "disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .hd_pmaif_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .pcs_rx_block_sel = "eightg";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .pcs_rx_clk_out_sel = "eightg_clk_out";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .pcs_rx_clk_sel = "pcs_rx_clk";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .pcs_rx_hip_clk_en = "hip_rx_disable";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .pcs_rx_output_sel = "teng_output";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_rx_pld_pcs_interface.inst_twentynm_hssi_rx_pld_pcs_interface .silicon_rev = "20nm5";

twentynm_hssi_common_pld_pcs_interface \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pldif_10g_rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
	.int_pldif_10g_tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
	.int_pldif_8g_rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
	.int_pldif_8g_tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
	.int_pldif_pmaif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
	.int_pldif_pmaif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
	.int_pldif_pmaif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
	.int_pldif_pmaif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
	.int_pldif_pmaif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
	.int_pldif_pmaif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
	.int_pldif_pmaif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
	.int_pldif_pmaif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
	.int_pldif_pmaif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
	.int_pldif_pmaif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
	.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
	.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
	.pld_8g_refclk_dig2(gnd),
	.pld_atpg_los_en_n(vcc),
	.pld_ltr(gnd),
	.pld_mem_krfec_atpg_rst_n(vcc),
	.pld_partial_reconfig(vcc),
	.pld_pcs_refclk_dig(gnd),
	.pld_pma_adapt_start(gnd),
	.pld_pma_csr_test_dis(vcc),
	.pld_pma_early_eios(gnd),
	.pld_pma_ltd_b(vcc),
	.pld_pma_nrpi_freeze(gnd),
	.pld_pma_ppm_lock(vcc),
	.pld_pma_rs_lpbk_b(!in_pld_pma_rs_lpbk_b),
	.pld_pma_rx_qpi_pullup(vcc),
	.pld_pma_tx_bitslip(gnd),
	.pld_pma_tx_bonding_rstb(gnd),
	.pld_pma_tx_qpi_pulldn(vcc),
	.pld_pma_tx_qpi_pullup(vcc),
	.pld_pma_txdetectrx(gnd),
	.pld_scan_mode_n(vcc),
	.pld_scan_shift_n(vcc),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.int_pldif_10g_test_data({\w_hssi_10g_tx_pcs_tx_test_data[19] ,\w_hssi_10g_tx_pcs_tx_test_data[18] ,\w_hssi_10g_tx_pcs_tx_test_data[17] ,\w_hssi_10g_tx_pcs_tx_test_data[16] ,\w_hssi_10g_tx_pcs_tx_test_data[15] ,\w_hssi_10g_tx_pcs_tx_test_data[14] ,\w_hssi_10g_tx_pcs_tx_test_data[13] ,
\w_hssi_10g_tx_pcs_tx_test_data[12] ,\w_hssi_10g_tx_pcs_tx_test_data[11] ,\w_hssi_10g_tx_pcs_tx_test_data[10] ,\w_hssi_10g_tx_pcs_tx_test_data[9] ,\w_hssi_10g_tx_pcs_tx_test_data[8] ,\w_hssi_10g_tx_pcs_tx_test_data[7] ,\w_hssi_10g_tx_pcs_tx_test_data[6] ,
\w_hssi_10g_tx_pcs_tx_test_data[5] ,\w_hssi_10g_tx_pcs_tx_test_data[4] ,\w_hssi_10g_tx_pcs_tx_test_data[3] ,\w_hssi_10g_tx_pcs_tx_test_data[2] ,\w_hssi_10g_tx_pcs_tx_test_data[1] ,\w_hssi_10g_tx_pcs_tx_test_data[0] }),
	.int_pldif_8g_chnl_test_bus_out({\w_hssi_8g_rx_pcs_chnl_test_bus_out[19] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[18] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[17] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[16] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[15] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[14] ,
\w_hssi_8g_rx_pcs_chnl_test_bus_out[13] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[12] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[11] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[10] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[9] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[8] ,
\w_hssi_8g_rx_pcs_chnl_test_bus_out[7] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[6] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[5] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[4] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[3] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[2] ,
\w_hssi_8g_rx_pcs_chnl_test_bus_out[1] ,\w_hssi_8g_rx_pcs_chnl_test_bus_out[0] }),
	.int_pldif_avmm_refclk_dig_en(),
	.int_pldif_g3_test_out({\w_hssi_pipe_gen3_test_out[19] ,\w_hssi_pipe_gen3_test_out[18] ,\w_hssi_pipe_gen3_test_out[17] ,\w_hssi_pipe_gen3_test_out[16] ,\w_hssi_pipe_gen3_test_out[15] ,\w_hssi_pipe_gen3_test_out[14] ,\w_hssi_pipe_gen3_test_out[13] ,\w_hssi_pipe_gen3_test_out[12] ,
\w_hssi_pipe_gen3_test_out[11] ,\w_hssi_pipe_gen3_test_out[10] ,\w_hssi_pipe_gen3_test_out[9] ,\w_hssi_pipe_gen3_test_out[8] ,\w_hssi_pipe_gen3_test_out[7] ,\w_hssi_pipe_gen3_test_out[6] ,\w_hssi_pipe_gen3_test_out[5] ,\w_hssi_pipe_gen3_test_out[4] ,
\w_hssi_pipe_gen3_test_out[3] ,\w_hssi_pipe_gen3_test_out[2] ,\w_hssi_pipe_gen3_test_out[1] ,\w_hssi_pipe_gen3_test_out[0] }),
	.int_pldif_krfec_test_data({\w_hssi_krfec_tx_pcs_tx_test_data[19] ,\w_hssi_krfec_tx_pcs_tx_test_data[18] ,\w_hssi_krfec_tx_pcs_tx_test_data[17] ,\w_hssi_krfec_tx_pcs_tx_test_data[16] ,\w_hssi_krfec_tx_pcs_tx_test_data[15] ,\w_hssi_krfec_tx_pcs_tx_test_data[14] ,
\w_hssi_krfec_tx_pcs_tx_test_data[13] ,\w_hssi_krfec_tx_pcs_tx_test_data[12] ,\w_hssi_krfec_tx_pcs_tx_test_data[11] ,\w_hssi_krfec_tx_pcs_tx_test_data[10] ,\w_hssi_krfec_tx_pcs_tx_test_data[9] ,\w_hssi_krfec_tx_pcs_tx_test_data[8] ,
\w_hssi_krfec_tx_pcs_tx_test_data[7] ,\w_hssi_krfec_tx_pcs_tx_test_data[6] ,\w_hssi_krfec_tx_pcs_tx_test_data[5] ,\w_hssi_krfec_tx_pcs_tx_test_data[4] ,\w_hssi_krfec_tx_pcs_tx_test_data[3] ,\w_hssi_krfec_tx_pcs_tx_test_data[2] ,
\w_hssi_krfec_tx_pcs_tx_test_data[1] ,\w_hssi_krfec_tx_pcs_tx_test_data[0] }),
	.int_pldif_pmaif_pcie_sw_done({\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[1] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pcie_sw_done[0] }),
	.int_pldif_pmaif_pma_reserved_in({\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[4] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[3] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[2] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[1] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_reserved_in[0] }),
	.int_pldif_pmaif_test_out({\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[19] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[18] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[17] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[16] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[15] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[14] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[13] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[12] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[11] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[10] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[9] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[8] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[7] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[6] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[5] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[4] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[3] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[2] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[1] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_test_out[0] }),
	.int_pldif_pmaif_testbus({\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[7] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[6] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[5] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[4] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[3] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[2] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[1] ,\w_hssi_common_pcs_pma_interface_int_pmaif_pldif_testbus[0] }),
	.pld_8g_eidleinfersel({gnd,gnd,gnd}),
	.pld_g3_current_coeff({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.pld_g3_current_rxpreset({gnd,gnd,gnd}),
	.pld_pma_eye_monitor({gnd,gnd,gnd,gnd,gnd,gnd}),
	.pld_pma_pcie_switch({gnd,gnd}),
	.pld_pma_reserved_out({vcc,gnd,gnd,gnd,gnd}),
	.pld_rate({gnd,gnd}),
	.pld_reserved_in({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.blockselect(out_blockselect_hssi_common_pld_pcs_interface),
	.hip_iocsr_rdy(),
	.hip_iocsr_rdy_dly(),
	.hip_nfrzdrv(),
	.hip_npor(),
	.hip_usermode(),
	.int_pldif_10g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
	.int_pldif_10g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
	.int_pldif_8g_ltr(),
	.int_pldif_8g_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
	.int_pldif_8g_refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
	.int_pldif_8g_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
	.int_pldif_avmm_pld_avmm1_request(),
	.int_pldif_avmm_pld_avmm2_request(),
	.int_pldif_g3_scan_mode_n(),
	.int_pldif_krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
	.int_pldif_krfec_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
	.int_pldif_krfec_scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
	.int_pldif_mem_atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
	.int_pldif_mem_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
	.int_pldif_pmaif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
	.int_pldif_pmaif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
	.int_pldif_pmaif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
	.int_pldif_pmaif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
	.int_pldif_pmaif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
	.int_pldif_pmaif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
	.int_pldif_pmaif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
	.int_pldif_pmaif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
	.int_pldif_pmaif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
	.int_pldif_pmaif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
	.int_pldif_pmaif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
	.int_pldif_pmaif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
	.int_pldif_pmaif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
	.int_pldif_pmaif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
	.int_pldif_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
	.int_pldif_pmaif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
	.int_pldif_pmaif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
	.int_pldif_pmaif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
	.int_pldif_pmaif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
	.int_pldif_pmaif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
	.int_pldif_pmaif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
	.int_pldif_pmaif_uhsif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
	.int_pldif_usr_rst_sel(w_hssi_common_pld_pcs_interface_int_pldif_usr_rst_sel),
	.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
	.pld_8g_eidleinfersel_fifo(),
	.pld_8g_eidleinfersel_reg(),
	.pld_partial_reconfig_fifo(),
	.pld_partial_reconfig_rx_div_by_2_rxclk_wire(),
	.pld_partial_reconfig_rx_div_by_2_txclk_wire(),
	.pld_partial_reconfig_rxclk_reg(),
	.pld_partial_reconfig_tx_div_by_2_wire(),
	.pld_partial_reconfig_txclk_reg(),
	.pld_pma_adapt_done(),
	.pld_pma_clklow(),
	.pld_pma_fref(),
	.pld_pma_hclk(),
	.pld_pma_pfdmode_lock(out_pld_pma_pfdmode_lock),
	.pld_pma_rx_detect_valid(),
	.pld_pma_rx_found(),
	.pld_pma_rxpll_lock(out_pld_pma_rxpll_lock),
	.pld_pmaif_mask_tx_pll(),
	.pld_rate_reg(),
	.pld_test_data_reg(),
	.pld_uhsif_lock(),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
	.avmmreaddata(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_AVMMREADDATA_bus ),
	.hip_cmn_clk(),
	.hip_cmn_ctrl(),
	.int_pldif_8g_eidleinfersel(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_8G_EIDLEINFERSEL_bus ),
	.int_pldif_g3_current_coeff(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_COEFF_bus ),
	.int_pldif_g3_current_rxpreset(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_G3_CURRENT_RXPRESET_bus ),
	.int_pldif_pmaif_eye_monitor(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_EYE_MONITOR_bus ),
	.int_pldif_pmaif_pcie_switch(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PCIE_SWITCH_bus ),
	.int_pldif_pmaif_pma_reserved_out(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_PMA_RESERVED_OUT_bus ),
	.int_pldif_pmaif_rate(\gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface_INT_PLDIF_PMAIF_RATE_bus ),
	.pld_pma_pcie_sw_done(),
	.pld_pma_reserved_in(),
	.pld_pma_testbus(),
	.pld_reserved_out(),
	.pld_test_data());
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .dft_clk_out_en = "dft_clk_out_disable";
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .dft_clk_out_sel = "teng_rx_dft_clk";
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .hrdrstctrl_en = "hrst_dis";
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .pcs_testbus_block_sel = "pma_if";
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_common_pld_pcs_interface.inst_twentynm_hssi_common_pld_pcs_interface .silicon_rev = "20nm5";

twentynm_hssi_tx_pld_pcs_interface \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pldif_10g_tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
	.int_pldif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
	.int_pldif_10g_tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
	.int_pldif_10g_tx_empty(w_hssi_10g_tx_pcs_tx_empty),
	.int_pldif_10g_tx_frame(w_hssi_10g_tx_pcs_tx_frame),
	.int_pldif_10g_tx_full(w_hssi_10g_tx_pcs_tx_full),
	.int_pldif_10g_tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
	.int_pldif_10g_tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
	.int_pldif_10g_tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
	.int_pldif_8g_empty_tx(w_hssi_8g_tx_pcs_ph_fifo_underflow),
	.int_pldif_8g_full_tx(w_hssi_8g_tx_pcs_ph_fifo_overflow),
	.int_pldif_8g_tx_clk_out(w_hssi_8g_tx_pcs_clk_out),
	.int_pldif_8g_tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
	.int_pldif_krfec_tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
	.int_pldif_krfec_tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
	.int_pldif_pmaif_clkdiv_tx(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
	.int_pldif_pmaif_clkdiv_tx_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
	.int_pldif_pmaif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
	.pld_10g_krfec_tx_pld_rst_n(!in_pld_10g_krfec_tx_pld_rst_n),
	.pld_10g_tx_burst_en(gnd),
	.pld_10g_tx_data_valid(gnd),
	.pld_10g_tx_wordslip(gnd),
	.pld_8g_g3_tx_pld_rst_n(!in_pld_10g_krfec_tx_pld_rst_n),
	.pld_8g_rddisable_tx(gnd),
	.pld_8g_wrenable_tx(gnd),
	.pld_partial_reconfig(vcc),
	.pld_pma_txpma_rstb(!in_pld_pma_txpma_rstb),
	.pld_pmaif_tx_pld_rst_n(!in_pld_10g_krfec_tx_pld_rst_n),
	.pld_polinv_tx(gnd),
	.pld_tx_clk(in_pld_tx_clk),
	.pld_txelecidle(gnd),
	.pld_uhsif_tx_clk(gnd),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_scan_mode_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.hip_tx_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.int_pldif_10g_tx_fifo_num({\w_hssi_10g_tx_pcs_tx_fifo_num[3] ,\w_hssi_10g_tx_pcs_tx_fifo_num[2] ,\w_hssi_10g_tx_pcs_tx_fifo_num[1] ,\w_hssi_10g_tx_pcs_tx_fifo_num[0] }),
	.pld_10g_tx_bitslip({gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.pld_10g_tx_diag_status({gnd,gnd}),
	.pld_8g_tx_boundary_sel({gnd,gnd,gnd,gnd,gnd}),
	.pld_tx_control({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.pld_tx_data({in_pld_tx_data[127],in_pld_tx_data[126],in_pld_tx_data[125],in_pld_tx_data[124],in_pld_tx_data[123],in_pld_tx_data[122],in_pld_tx_data[121],in_pld_tx_data[120],in_pld_tx_data[119],in_pld_tx_data[118],in_pld_tx_data[117],in_pld_tx_data[116],in_pld_tx_data[115],in_pld_tx_data[114],in_pld_tx_data[113],in_pld_tx_data[112],in_pld_tx_data[111],in_pld_tx_data[110],
in_pld_tx_data[109],in_pld_tx_data[108],in_pld_tx_data[107],in_pld_tx_data[106],in_pld_tx_data[105],in_pld_tx_data[104],in_pld_tx_data[103],in_pld_tx_data[102],in_pld_tx_data[101],in_pld_tx_data[100],in_pld_tx_data[99],in_pld_tx_data[98],in_pld_tx_data[97],in_pld_tx_data[96],in_pld_tx_data[95],in_pld_tx_data[94],in_pld_tx_data[93],in_pld_tx_data[92],
in_pld_tx_data[91],in_pld_tx_data[90],in_pld_tx_data[89],in_pld_tx_data[88],in_pld_tx_data[87],in_pld_tx_data[86],in_pld_tx_data[85],in_pld_tx_data[84],in_pld_tx_data[83],in_pld_tx_data[82],in_pld_tx_data[81],in_pld_tx_data[80],in_pld_tx_data[79],in_pld_tx_data[78],in_pld_tx_data[77],in_pld_tx_data[76],in_pld_tx_data[75],in_pld_tx_data[74],
in_pld_tx_data[73],in_pld_tx_data[72],in_pld_tx_data[71],in_pld_tx_data[70],in_pld_tx_data[69],in_pld_tx_data[68],in_pld_tx_data[67],in_pld_tx_data[66],in_pld_tx_data[65],in_pld_tx_data[64],in_pld_tx_data[63],in_pld_tx_data[62],in_pld_tx_data[61],in_pld_tx_data[60],in_pld_tx_data[59],in_pld_tx_data[58],in_pld_tx_data[57],in_pld_tx_data[56],
in_pld_tx_data[55],in_pld_tx_data[54],in_pld_tx_data[53],in_pld_tx_data[52],in_pld_tx_data[51],in_pld_tx_data[50],in_pld_tx_data[49],in_pld_tx_data[48],in_pld_tx_data[47],in_pld_tx_data[46],in_pld_tx_data[45],in_pld_tx_data[44],in_pld_tx_data[43],in_pld_tx_data[42],in_pld_tx_data[41],in_pld_tx_data[40],in_pld_tx_data[39],in_pld_tx_data[38],
in_pld_tx_data[37],in_pld_tx_data[36],in_pld_tx_data[35],in_pld_tx_data[34],in_pld_tx_data[33],in_pld_tx_data[32],in_pld_tx_data[31],in_pld_tx_data[30],in_pld_tx_data[29],in_pld_tx_data[28],in_pld_tx_data[27],in_pld_tx_data[26],in_pld_tx_data[25],in_pld_tx_data[24],in_pld_tx_data[23],in_pld_tx_data[22],in_pld_tx_data[21],in_pld_tx_data[20],
in_pld_tx_data[19],in_pld_tx_data[18],in_pld_tx_data[17],in_pld_tx_data[16],in_pld_tx_data[15],in_pld_tx_data[14],in_pld_tx_data[13],in_pld_tx_data[12],in_pld_tx_data[11],in_pld_tx_data[10],in_pld_tx_data[9],in_pld_tx_data[8],in_pld_tx_data[7],in_pld_tx_data[6],in_pld_tx_data[5],in_pld_tx_data[4],in_pld_tx_data[3],in_pld_tx_data[2],
in_pld_tx_data[1],in_pld_tx_data[0]}),
	.blockselect(out_blockselect_hssi_tx_pld_pcs_interface),
	.hip_clk_out_div_by_2_wire(),
	.hip_clk_out_wire(),
	.hip_tx_clk(),
	.int_pldif_10g_tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
	.int_pldif_10g_tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
	.int_pldif_10g_tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
	.int_pldif_10g_tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
	.int_pldif_10g_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
	.int_pldif_10g_tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
	.int_pldif_8g_pld_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
	.int_pldif_8g_rddisable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
	.int_pldif_8g_rev_loopbk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
	.int_pldif_8g_txdeemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
	.int_pldif_8g_txdetectrxloopback(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
	.int_pldif_8g_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
	.int_pldif_8g_txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
	.int_pldif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
	.int_pldif_8g_wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
	.int_pldif_pmaif_8g_txurstpcs_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
	.int_pldif_pmaif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
	.int_pldif_pmaif_tx_pld_clk(),
	.int_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
	.int_pldif_pmaif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
	.int_pldif_pmaif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
	.int_pldif_pmaif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
	.pld_10g_krfec_tx_frame(),
	.pld_10g_tx_burst_en_exe(),
	.pld_10g_tx_burst_en_exe_10g_fastreg(),
	.pld_10g_tx_burst_en_exe_plddirect_reg(),
	.pld_10g_tx_data_valid_2ff_delay1_fastreg(),
	.pld_10g_tx_data_valid_2ff_delay3_fastreg(),
	.pld_10g_tx_data_valid_2ff_delay4_fastreg(),
	.pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg(),
	.pld_10g_tx_data_valid_2ff_delay6_fastreg(),
	.pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg(),
	.pld_10g_tx_data_valid_fastreg(),
	.pld_10g_tx_data_valid_plddirect_fastreg(),
	.pld_10g_tx_empty(),
	.pld_10g_tx_full(),
	.pld_10g_tx_pempty(),
	.pld_10g_tx_pfull(),
	.pld_10g_tx_wordslip_exe(),
	.pld_8g_empty_tx(),
	.pld_8g_full_tx(),
	.pld_krfec_tx_alignment(),
	.pld_pcs_tx_clk_out(out_pld_pcs_tx_clk_out),
	.pld_pcs_tx_clk_out_pma_wire(),
	.pld_pma_clkdiv_tx_user(),
	.pld_pma_tx_clk_out(),
	.pld_pma_tx_clk_out_wire(),
	.pld_pmaif_tx_pld_rst_n_reg(),
	.pld_polinv_tx_10g_pcsdirect_reg(),
	.pld_polinv_tx_8g_reg(),
	.pld_polinv_tx_pat_reg(),
	.pld_tx_clk_fifo(),
	.pld_tx_control_fifo(),
	.pld_tx_control_hi_10g_reg(),
	.pld_tx_control_lo_10g_2ff_delay4_fastreg(),
	.pld_tx_control_lo_10g_2ff_delay6_fastreg(),
	.pld_tx_control_lo_10g_fastreg(),
	.pld_tx_control_lo_8g_2ff_delay4_fastreg(),
	.pld_tx_control_lo_8g_2ff_delay6_fastreg(),
	.pld_tx_control_lo_8g_fastreg(),
	.pld_tx_control_lo_plddirect_2ff_delay1_fastreg(),
	.pld_tx_control_lo_plddirect_2ff_delay3_fastreg(),
	.pld_tx_control_lo_plddirect_2ff_delay4_fastreg(),
	.pld_tx_control_lo_plddirect_2ff_delay6_fastreg(),
	.pld_tx_control_lo_plddirect_fastreg(),
	.pld_tx_control_lo_plddirect_reg(),
	.pld_tx_data_hi_reg(),
	.pld_tx_data_lo_10g_2ff_delay4_fastreg(),
	.pld_tx_data_lo_10g_2ff_delay6_fastreg(),
	.pld_tx_data_lo_10g_fastreg(),
	.pld_tx_data_lo_8g_2ff_delay4_fastreg(),
	.pld_tx_data_lo_8g_2ff_delay6_fastreg(),
	.pld_tx_data_lo_8g_fastreg(),
	.pld_tx_data_lo_plddirect_2ff_delay1_fastreg(),
	.pld_tx_data_lo_plddirect_2ff_delay3_fastreg(),
	.pld_tx_data_lo_plddirect_2ff_delay4_fastreg(),
	.pld_tx_data_lo_plddirect_2ff_delay6_fastreg(),
	.pld_tx_data_lo_plddirect_fastreg(),
	.pld_tx_data_lo_plddirect_reg(),
	.pld_uhsif_reg(),
	.pld_uhsif_tx_clk_out(),
	.pma_tx_pma_clk_reg(),
	.avmmreaddata(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_AVMMREADDATA_bus ),
	.int_pldif_10g_tx_bitslip(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_BITSLIP_bus ),
	.int_pldif_10g_tx_control(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_bus ),
	.int_pldif_10g_tx_control_reg(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_CONTROL_REG_bus ),
	.int_pldif_10g_tx_data(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_bus ),
	.int_pldif_10g_tx_data_reg(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DATA_REG_bus ),
	.int_pldif_10g_tx_diag_status(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_10G_TX_DIAG_STATUS_bus ),
	.int_pldif_8g_powerdown(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_POWERDOWN_bus ),
	.int_pldif_8g_tx_blk_start(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BLK_START_bus ),
	.int_pldif_8g_tx_boundary_sel(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_BOUNDARY_SEL_bus ),
	.int_pldif_8g_tx_data_valid(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_DATA_VALID_bus ),
	.int_pldif_8g_tx_sync_hdr(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TX_SYNC_HDR_bus ),
	.int_pldif_8g_txd(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_bus ),
	.int_pldif_8g_txd_fast_reg(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXD_FAST_REG_bus ),
	.int_pldif_8g_txmargin(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_8G_TXMARGIN_bus ),
	.int_pldif_pmaif_tx_data(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_TX_DATA_bus ),
	.int_pldif_pmaif_uhsif_tx_data(\gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface_INT_PLDIF_PMAIF_UHSIF_TX_DATA_bus ),
	.pld_10g_tx_fifo_num());
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_advanced_user_mode_tx = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_ctrl_plane_bonding_tx = "individual_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_fifo_mode_tx = "fifo_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_low_latency_en_tx = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_pma_dw_tx = "pma_64b_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_prot_mode_tx = "disabled_prot_mode_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_shared_fifo_width_tx = "single_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_10g_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_ctrl_plane_bonding_tx = "individual_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_fifo_mode_tx = "reg_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_hip_mode = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_pma_dw_tx = "pma_10b_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_prot_mode_tx = "cpri_rx_tx_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_8g_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_ctrl_plane_bonding_tx = "individual_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_frequency_rules_en = "enable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_func_mode = "enable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_hclk_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_hip_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_hrdrstctl_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_low_latency_en_tx = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pcs_tx_ac_pwr_uw_per_mhz = 20'b00000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pcs_tx_pwr_scaling_clk = "pma_tx_clk";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pld_fifo_mode_tx = "reg_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pld_tx_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pld_uhsif_tx_clk_hz = 30'b000000000000000000000000000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pma_dw_tx = "pma_10b_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_pma_tx_clk_hz = 30'b000111011100110101100101000000;
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_prot_mode_tx = "cpri_8b10b_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_shared_fifo_width_tx = "single_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_speed_grade = "e2";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_chnl_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_fifo_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_fifo_prot_mode_tx = "non_teng_mode_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_fifo_shared_fifo_width_tx = "single_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_fifo_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_g3_prot_mode = "disabled_prot_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_g3_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_krfec_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_krfec_low_latency_en_tx = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_krfec_lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_krfec_prot_mode_tx = "disabled_prot_mode_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_krfec_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pldif_hrdrstctl_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pldif_prot_mode_tx = "eightg_and_g3_reg_mode_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pldif_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_ctrl_plane_bonding = "individual";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_pma_dw_tx = "pma_10b_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_prot_mode_tx = "eightg_only_pld_mode_tx";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_sim_mode = "disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .hd_pmaif_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_clk_out_sel = "eightg_clk_out";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_clk_source = "eightg";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_data_source = "hip_disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay1_clk_en = "delay1_clk_disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay1_clk_sel = "pcs_tx_clk";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay1_ctrl = "delay1_path0";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay1_data_sel = "one_ff_delay";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay2_clk_en = "delay2_clk_disable";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_delay2_ctrl = "delay2_path0";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .pcs_tx_output_sel = "teng_output";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_tx_pld_pcs_interface.inst_twentynm_hssi_tx_pld_pcs_interface .silicon_rev = "20nm5";

twentynm_hssi_10g_rx_pcs \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
	.rx_align_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_align_clr),
	.rx_bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_bitslip),
	.rx_clr_ber_count(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_ber_count),
	.rx_clr_errblk_cnt(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_clr_errblk_cnt),
	.rx_data_valid_fb(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_valid_fb),
	.rx_data_valid_in_krfec(w_hssi_krfec_rx_pcs_rx_data_valid_out),
	.rx_pld_clk(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_clk),
	.rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_pld_rst_n),
	.rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
	.rx_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_prbs_err_clr),
	.rx_rd_en(w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_rd_en),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
	.signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
	.signal_ok_krfec(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
	.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.r_rx_diag_word({gnd,vcc,vcc,gnd,gnd,vcc,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.r_rx_scrm_word({gnd,gnd,vcc,gnd,vcc,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.r_rx_skip_word({gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd}),
	.r_rx_sync_word({gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd}),
	.rx_control_fb({\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[19] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[18] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[17] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[16] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[15] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[14] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[13] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[12] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[11] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[10] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[9] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[8] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[7] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[6] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[5] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[4] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[3] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[2] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[1] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_control_fb[0] }),
	.rx_control_in_krfec({\w_hssi_krfec_rx_pcs_rx_control_out[9] ,\w_hssi_krfec_rx_pcs_rx_control_out[8] ,\w_hssi_krfec_rx_pcs_rx_control_out[7] ,\w_hssi_krfec_rx_pcs_rx_control_out[6] ,\w_hssi_krfec_rx_pcs_rx_control_out[5] ,\w_hssi_krfec_rx_pcs_rx_control_out[4] ,
\w_hssi_krfec_rx_pcs_rx_control_out[3] ,\w_hssi_krfec_rx_pcs_rx_control_out[2] ,\w_hssi_krfec_rx_pcs_rx_control_out[1] ,\w_hssi_krfec_rx_pcs_rx_control_out[0] }),
	.rx_data_fb({\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[127] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[126] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[125] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[124] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[123] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[122] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[121] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[120] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[119] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[118] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[117] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[116] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[115] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[114] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[113] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[112] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[111] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[110] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[109] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[108] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[107] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[106] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[105] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[104] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[103] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[102] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[101] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[100] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[99] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[98] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[97] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[96] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[95] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[94] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[93] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[92] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[91] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[90] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[89] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[88] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[87] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[86] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[85] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[84] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[83] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[82] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[81] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[80] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[79] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[78] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[77] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[76] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[75] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[74] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[73] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[72] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[71] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[70] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[69] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[68] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[67] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[66] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[65] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[64] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[63] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[62] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[61] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[60] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[59] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[58] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[57] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[56] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[55] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[54] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[53] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[52] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[51] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[50] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[49] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[48] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[47] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[46] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[45] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[44] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[43] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[42] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[41] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[40] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[39] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[38] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[37] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[36] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[35] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[34] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[33] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[32] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[31] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[30] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[29] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[28] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[27] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[26] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[25] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[24] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[23] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[22] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[21] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[20] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[19] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[18] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[17] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[16] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[15] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[14] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[13] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[12] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[11] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[10] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[9] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[8] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[7] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[6] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[5] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[4] ,
\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[3] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[2] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[1] ,\w_hssi_rx_pld_pcs_interface_int_pldif_10g_rx_data_fb[0] }),
	.rx_data_in_krfec({\w_hssi_krfec_rx_pcs_rx_data_out[63] ,\w_hssi_krfec_rx_pcs_rx_data_out[62] ,\w_hssi_krfec_rx_pcs_rx_data_out[61] ,\w_hssi_krfec_rx_pcs_rx_data_out[60] ,\w_hssi_krfec_rx_pcs_rx_data_out[59] ,\w_hssi_krfec_rx_pcs_rx_data_out[58] ,
\w_hssi_krfec_rx_pcs_rx_data_out[57] ,\w_hssi_krfec_rx_pcs_rx_data_out[56] ,\w_hssi_krfec_rx_pcs_rx_data_out[55] ,\w_hssi_krfec_rx_pcs_rx_data_out[54] ,\w_hssi_krfec_rx_pcs_rx_data_out[53] ,\w_hssi_krfec_rx_pcs_rx_data_out[52] ,
\w_hssi_krfec_rx_pcs_rx_data_out[51] ,\w_hssi_krfec_rx_pcs_rx_data_out[50] ,\w_hssi_krfec_rx_pcs_rx_data_out[49] ,\w_hssi_krfec_rx_pcs_rx_data_out[48] ,\w_hssi_krfec_rx_pcs_rx_data_out[47] ,\w_hssi_krfec_rx_pcs_rx_data_out[46] ,
\w_hssi_krfec_rx_pcs_rx_data_out[45] ,\w_hssi_krfec_rx_pcs_rx_data_out[44] ,\w_hssi_krfec_rx_pcs_rx_data_out[43] ,\w_hssi_krfec_rx_pcs_rx_data_out[42] ,\w_hssi_krfec_rx_pcs_rx_data_out[41] ,\w_hssi_krfec_rx_pcs_rx_data_out[40] ,
\w_hssi_krfec_rx_pcs_rx_data_out[39] ,\w_hssi_krfec_rx_pcs_rx_data_out[38] ,\w_hssi_krfec_rx_pcs_rx_data_out[37] ,\w_hssi_krfec_rx_pcs_rx_data_out[36] ,\w_hssi_krfec_rx_pcs_rx_data_out[35] ,\w_hssi_krfec_rx_pcs_rx_data_out[34] ,
\w_hssi_krfec_rx_pcs_rx_data_out[33] ,\w_hssi_krfec_rx_pcs_rx_data_out[32] ,\w_hssi_krfec_rx_pcs_rx_data_out[31] ,\w_hssi_krfec_rx_pcs_rx_data_out[30] ,\w_hssi_krfec_rx_pcs_rx_data_out[29] ,\w_hssi_krfec_rx_pcs_rx_data_out[28] ,
\w_hssi_krfec_rx_pcs_rx_data_out[27] ,\w_hssi_krfec_rx_pcs_rx_data_out[26] ,\w_hssi_krfec_rx_pcs_rx_data_out[25] ,\w_hssi_krfec_rx_pcs_rx_data_out[24] ,\w_hssi_krfec_rx_pcs_rx_data_out[23] ,\w_hssi_krfec_rx_pcs_rx_data_out[22] ,
\w_hssi_krfec_rx_pcs_rx_data_out[21] ,\w_hssi_krfec_rx_pcs_rx_data_out[20] ,\w_hssi_krfec_rx_pcs_rx_data_out[19] ,\w_hssi_krfec_rx_pcs_rx_data_out[18] ,\w_hssi_krfec_rx_pcs_rx_data_out[17] ,\w_hssi_krfec_rx_pcs_rx_data_out[16] ,
\w_hssi_krfec_rx_pcs_rx_data_out[15] ,\w_hssi_krfec_rx_pcs_rx_data_out[14] ,\w_hssi_krfec_rx_pcs_rx_data_out[13] ,\w_hssi_krfec_rx_pcs_rx_data_out[12] ,\w_hssi_krfec_rx_pcs_rx_data_out[11] ,\w_hssi_krfec_rx_pcs_rx_data_out[10] ,
\w_hssi_krfec_rx_pcs_rx_data_out[9] ,\w_hssi_krfec_rx_pcs_rx_data_out[8] ,\w_hssi_krfec_rx_pcs_rx_data_out[7] ,\w_hssi_krfec_rx_pcs_rx_data_out[6] ,\w_hssi_krfec_rx_pcs_rx_data_out[5] ,\w_hssi_krfec_rx_pcs_rx_data_out[4] ,\w_hssi_krfec_rx_pcs_rx_data_out[3] ,
\w_hssi_krfec_rx_pcs_rx_data_out[2] ,\w_hssi_krfec_rx_pcs_rx_data_out[1] ,\w_hssi_krfec_rx_pcs_rx_data_out[0] }),
	.rx_fifo_rd_data({\w_hssi_fifo_rx_pcs_data_out_10g[73] ,\w_hssi_fifo_rx_pcs_data_out_10g[72] ,\w_hssi_fifo_rx_pcs_data_out_10g[71] ,\w_hssi_fifo_rx_pcs_data_out_10g[70] ,\w_hssi_fifo_rx_pcs_data_out_10g[69] ,\w_hssi_fifo_rx_pcs_data_out_10g[68] ,
\w_hssi_fifo_rx_pcs_data_out_10g[67] ,\w_hssi_fifo_rx_pcs_data_out_10g[66] ,\w_hssi_fifo_rx_pcs_data_out_10g[65] ,\w_hssi_fifo_rx_pcs_data_out_10g[64] ,\w_hssi_fifo_rx_pcs_data_out_10g[63] ,\w_hssi_fifo_rx_pcs_data_out_10g[62] ,
\w_hssi_fifo_rx_pcs_data_out_10g[61] ,\w_hssi_fifo_rx_pcs_data_out_10g[60] ,\w_hssi_fifo_rx_pcs_data_out_10g[59] ,\w_hssi_fifo_rx_pcs_data_out_10g[58] ,\w_hssi_fifo_rx_pcs_data_out_10g[57] ,\w_hssi_fifo_rx_pcs_data_out_10g[56] ,
\w_hssi_fifo_rx_pcs_data_out_10g[55] ,\w_hssi_fifo_rx_pcs_data_out_10g[54] ,\w_hssi_fifo_rx_pcs_data_out_10g[53] ,\w_hssi_fifo_rx_pcs_data_out_10g[52] ,\w_hssi_fifo_rx_pcs_data_out_10g[51] ,\w_hssi_fifo_rx_pcs_data_out_10g[50] ,
\w_hssi_fifo_rx_pcs_data_out_10g[49] ,\w_hssi_fifo_rx_pcs_data_out_10g[48] ,\w_hssi_fifo_rx_pcs_data_out_10g[47] ,\w_hssi_fifo_rx_pcs_data_out_10g[46] ,\w_hssi_fifo_rx_pcs_data_out_10g[45] ,\w_hssi_fifo_rx_pcs_data_out_10g[44] ,
\w_hssi_fifo_rx_pcs_data_out_10g[43] ,\w_hssi_fifo_rx_pcs_data_out_10g[42] ,\w_hssi_fifo_rx_pcs_data_out_10g[41] ,\w_hssi_fifo_rx_pcs_data_out_10g[40] ,\w_hssi_fifo_rx_pcs_data_out_10g[39] ,\w_hssi_fifo_rx_pcs_data_out_10g[38] ,
\w_hssi_fifo_rx_pcs_data_out_10g[37] ,\w_hssi_fifo_rx_pcs_data_out_10g[36] ,\w_hssi_fifo_rx_pcs_data_out_10g[35] ,\w_hssi_fifo_rx_pcs_data_out_10g[34] ,\w_hssi_fifo_rx_pcs_data_out_10g[33] ,\w_hssi_fifo_rx_pcs_data_out_10g[32] ,
\w_hssi_fifo_rx_pcs_data_out_10g[31] ,\w_hssi_fifo_rx_pcs_data_out_10g[30] ,\w_hssi_fifo_rx_pcs_data_out_10g[29] ,\w_hssi_fifo_rx_pcs_data_out_10g[28] ,\w_hssi_fifo_rx_pcs_data_out_10g[27] ,\w_hssi_fifo_rx_pcs_data_out_10g[26] ,
\w_hssi_fifo_rx_pcs_data_out_10g[25] ,\w_hssi_fifo_rx_pcs_data_out_10g[24] ,\w_hssi_fifo_rx_pcs_data_out_10g[23] ,\w_hssi_fifo_rx_pcs_data_out_10g[22] ,\w_hssi_fifo_rx_pcs_data_out_10g[21] ,\w_hssi_fifo_rx_pcs_data_out_10g[20] ,
\w_hssi_fifo_rx_pcs_data_out_10g[19] ,\w_hssi_fifo_rx_pcs_data_out_10g[18] ,\w_hssi_fifo_rx_pcs_data_out_10g[17] ,\w_hssi_fifo_rx_pcs_data_out_10g[16] ,\w_hssi_fifo_rx_pcs_data_out_10g[15] ,\w_hssi_fifo_rx_pcs_data_out_10g[14] ,
\w_hssi_fifo_rx_pcs_data_out_10g[13] ,\w_hssi_fifo_rx_pcs_data_out_10g[12] ,\w_hssi_fifo_rx_pcs_data_out_10g[11] ,\w_hssi_fifo_rx_pcs_data_out_10g[10] ,\w_hssi_fifo_rx_pcs_data_out_10g[9] ,\w_hssi_fifo_rx_pcs_data_out_10g[8] ,\w_hssi_fifo_rx_pcs_data_out_10g[7] ,
\w_hssi_fifo_rx_pcs_data_out_10g[6] ,\w_hssi_fifo_rx_pcs_data_out_10g[5] ,\w_hssi_fifo_rx_pcs_data_out_10g[4] ,\w_hssi_fifo_rx_pcs_data_out_10g[3] ,\w_hssi_fifo_rx_pcs_data_out_10g[2] ,\w_hssi_fifo_rx_pcs_data_out_10g[1] ,\w_hssi_fifo_rx_pcs_data_out_10g[0] }),
	.rx_fifo_rd_data_dw({\w_hssi_fifo_rx_pcs_data_out2_10g[73] ,\w_hssi_fifo_rx_pcs_data_out2_10g[72] ,\w_hssi_fifo_rx_pcs_data_out2_10g[71] ,\w_hssi_fifo_rx_pcs_data_out2_10g[70] ,\w_hssi_fifo_rx_pcs_data_out2_10g[69] ,\w_hssi_fifo_rx_pcs_data_out2_10g[68] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[67] ,\w_hssi_fifo_rx_pcs_data_out2_10g[66] ,\w_hssi_fifo_rx_pcs_data_out2_10g[65] ,\w_hssi_fifo_rx_pcs_data_out2_10g[64] ,\w_hssi_fifo_rx_pcs_data_out2_10g[63] ,\w_hssi_fifo_rx_pcs_data_out2_10g[62] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[61] ,\w_hssi_fifo_rx_pcs_data_out2_10g[60] ,\w_hssi_fifo_rx_pcs_data_out2_10g[59] ,\w_hssi_fifo_rx_pcs_data_out2_10g[58] ,\w_hssi_fifo_rx_pcs_data_out2_10g[57] ,\w_hssi_fifo_rx_pcs_data_out2_10g[56] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[55] ,\w_hssi_fifo_rx_pcs_data_out2_10g[54] ,\w_hssi_fifo_rx_pcs_data_out2_10g[53] ,\w_hssi_fifo_rx_pcs_data_out2_10g[52] ,\w_hssi_fifo_rx_pcs_data_out2_10g[51] ,\w_hssi_fifo_rx_pcs_data_out2_10g[50] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[49] ,\w_hssi_fifo_rx_pcs_data_out2_10g[48] ,\w_hssi_fifo_rx_pcs_data_out2_10g[47] ,\w_hssi_fifo_rx_pcs_data_out2_10g[46] ,\w_hssi_fifo_rx_pcs_data_out2_10g[45] ,\w_hssi_fifo_rx_pcs_data_out2_10g[44] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[43] ,\w_hssi_fifo_rx_pcs_data_out2_10g[42] ,\w_hssi_fifo_rx_pcs_data_out2_10g[41] ,\w_hssi_fifo_rx_pcs_data_out2_10g[40] ,\w_hssi_fifo_rx_pcs_data_out2_10g[39] ,\w_hssi_fifo_rx_pcs_data_out2_10g[38] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[37] ,\w_hssi_fifo_rx_pcs_data_out2_10g[36] ,\w_hssi_fifo_rx_pcs_data_out2_10g[35] ,\w_hssi_fifo_rx_pcs_data_out2_10g[34] ,\w_hssi_fifo_rx_pcs_data_out2_10g[33] ,\w_hssi_fifo_rx_pcs_data_out2_10g[32] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[31] ,\w_hssi_fifo_rx_pcs_data_out2_10g[30] ,\w_hssi_fifo_rx_pcs_data_out2_10g[29] ,\w_hssi_fifo_rx_pcs_data_out2_10g[28] ,\w_hssi_fifo_rx_pcs_data_out2_10g[27] ,\w_hssi_fifo_rx_pcs_data_out2_10g[26] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[25] ,\w_hssi_fifo_rx_pcs_data_out2_10g[24] ,\w_hssi_fifo_rx_pcs_data_out2_10g[23] ,\w_hssi_fifo_rx_pcs_data_out2_10g[22] ,\w_hssi_fifo_rx_pcs_data_out2_10g[21] ,\w_hssi_fifo_rx_pcs_data_out2_10g[20] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[19] ,\w_hssi_fifo_rx_pcs_data_out2_10g[18] ,\w_hssi_fifo_rx_pcs_data_out2_10g[17] ,\w_hssi_fifo_rx_pcs_data_out2_10g[16] ,\w_hssi_fifo_rx_pcs_data_out2_10g[15] ,\w_hssi_fifo_rx_pcs_data_out2_10g[14] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[13] ,\w_hssi_fifo_rx_pcs_data_out2_10g[12] ,\w_hssi_fifo_rx_pcs_data_out2_10g[11] ,\w_hssi_fifo_rx_pcs_data_out2_10g[10] ,\w_hssi_fifo_rx_pcs_data_out2_10g[9] ,\w_hssi_fifo_rx_pcs_data_out2_10g[8] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[7] ,\w_hssi_fifo_rx_pcs_data_out2_10g[6] ,\w_hssi_fifo_rx_pcs_data_out2_10g[5] ,\w_hssi_fifo_rx_pcs_data_out2_10g[4] ,\w_hssi_fifo_rx_pcs_data_out2_10g[3] ,\w_hssi_fifo_rx_pcs_data_out2_10g[2] ,
\w_hssi_fifo_rx_pcs_data_out2_10g[1] ,\w_hssi_fifo_rx_pcs_data_out2_10g[0] }),
	.rx_pma_data({\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[63] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[62] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[61] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[60] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[59] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[58] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[57] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[56] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[55] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[54] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[53] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[52] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[51] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[50] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[49] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[48] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[47] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[46] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[45] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[44] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[43] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[42] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[41] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[40] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[39] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[38] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[37] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[36] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[35] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[34] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[33] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[32] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[31] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[30] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[29] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[28] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[27] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[26] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[25] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[24] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[23] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[22] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[21] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[20] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[19] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[18] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[17] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[16] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[15] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[14] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[13] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[12] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[11] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[10] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[9] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[8] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[7] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[6] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[5] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[4] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[3] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[2] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[1] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_data[0] }),
	.blockselect(out_blockselect_hssi_10g_rx_pcs),
	.pld_10g_krfec_rx_blk_lock_10g_reg(),
	.pld_10g_krfec_rx_blk_lock_10g_txclk_reg(),
	.pld_10g_krfec_rx_clr_errblk_cnt_reg(),
	.pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg(),
	.pld_10g_krfec_rx_diag_data_status_10g_reg(),
	.pld_10g_krfec_rx_diag_data_status_10g_txclk_reg(),
	.pld_10g_krfec_rx_frame_10g_reg(),
	.pld_10g_krfec_rx_frame_10g_txclk_reg(),
	.pld_10g_krfec_rx_pld_rst_n_fifo(),
	.pld_10g_krfec_rx_pld_rst_n_reg(),
	.pld_10g_krfec_rx_pld_rst_n_txclk_reg(),
	.pld_10g_rx_align_clr_fifo(),
	.pld_10g_rx_align_clr_reg(),
	.pld_10g_rx_align_clr_txclk_reg(),
	.pld_10g_rx_align_val_fifo(),
	.pld_10g_rx_align_val_reg(),
	.pld_10g_rx_align_val_txclk_reg(),
	.pld_10g_rx_clr_ber_count_reg(),
	.pld_10g_rx_clr_ber_count_txclk_reg(),
	.pld_10g_rx_crc32_err_reg(),
	.pld_10g_rx_crc32_err_txclk_reg(),
	.pld_10g_rx_data_valid_10g_reg(),
	.pld_10g_rx_data_valid_fifo(),
	.pld_10g_rx_data_valid_pcsdirect_reg(),
	.pld_10g_rx_data_valid_txclk_reg(),
	.pld_10g_rx_empty_fifo(),
	.pld_10g_rx_fifo_del_reg(),
	.pld_10g_rx_fifo_del_txclk_reg(),
	.pld_10g_rx_fifo_insert_fifo(),
	.pld_10g_rx_fifo_num_reg(),
	.pld_10g_rx_fifo_num_txclk_reg(),
	.pld_10g_rx_frame_lock_reg(),
	.pld_10g_rx_frame_lock_txclk_reg(),
	.pld_10g_rx_hi_ber_reg(),
	.pld_10g_rx_hi_ber_txclk_reg(),
	.pld_10g_rx_oflw_err_reg(),
	.pld_10g_rx_oflw_err_txclk_reg(),
	.pld_10g_rx_pempty_fifo(),
	.pld_10g_rx_pfull_reg(),
	.pld_10g_rx_pfull_txclk_reg(),
	.pld_10g_rx_rd_en_fifo(),
	.pld_pcs_rx_clk_out_10g_txclk_wire(),
	.pld_pcs_rx_clk_out_10g_wire(),
	.pld_rx_control_10g_reg(),
	.pld_rx_control_10g_txclk_reg(),
	.pld_rx_data_10g_reg(),
	.pld_rx_data_10g_txclk_reg(),
	.pld_rx_prbs_err_10g_txclk_reg(),
	.pld_rx_prbs_err_clr_10g_txclk_reg(),
	.rx_align_val(w_hssi_10g_rx_pcs_rx_align_val),
	.rx_blk_lock(w_hssi_10g_rx_pcs_rx_blk_lock),
	.rx_clk_out(w_hssi_10g_rx_pcs_rx_clk_out),
	.rx_clk_out_pld_if(w_hssi_10g_rx_pcs_rx_clk_out_pld_if),
	.rx_crc32_err(w_hssi_10g_rx_pcs_rx_crc32_err),
	.rx_data_valid(w_hssi_10g_rx_pcs_rx_data_valid),
	.rx_dft_clk_out(w_hssi_10g_rx_pcs_rx_dft_clk_out),
	.rx_empty(w_hssi_10g_rx_pcs_rx_empty),
	.rx_fec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
	.rx_fifo_del(w_hssi_10g_rx_pcs_rx_fifo_del),
	.rx_fifo_insert(w_hssi_10g_rx_pcs_rx_fifo_insert),
	.rx_fifo_wr_clk(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
	.rx_fifo_wr_en(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
	.rx_fifo_wr_rst_n(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
	.rx_frame_lock(w_hssi_10g_rx_pcs_rx_frame_lock),
	.rx_hi_ber(w_hssi_10g_rx_pcs_rx_hi_ber),
	.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
	.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
	.rx_oflw_err(w_hssi_10g_rx_pcs_rx_oflw_err),
	.rx_pempty(w_hssi_10g_rx_pcs_rx_pempty),
	.rx_pfull(w_hssi_10g_rx_pcs_rx_pfull),
	.rx_random_err(w_hssi_10g_rx_pcs_rx_random_err),
	.rx_rx_frame(w_hssi_10g_rx_pcs_rx_rx_frame),
	.avmmreaddata(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_AVMMREADDATA_bus ),
	.rx_control(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_CONTROL_bus ),
	.rx_data(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DATA_bus ),
	.rx_diag_status(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_DIAG_STATUS_bus ),
	.rx_fifo_num(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_NUM_bus ),
	.rx_fifo_rd_ptr(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR_bus ),
	.rx_fifo_rd_ptr2(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_RD_PTR2_bus ),
	.rx_fifo_wr_data(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_DATA_bus ),
	.rx_fifo_wr_ptr(\gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs_RX_FIFO_WR_PTR_bus ),
	.rx_test_data());
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .advanced_user_mode = "disable";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .align_del = "align_del_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .ber_bit_err_total_cnt = "bit_err_total_cnt_10g";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .ber_clken = "ber_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .ber_xus_timer_window = 21'b000000100110001001010;
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .bitslip_mode = "bitslip_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_bitslip_type = "bitslip_comb";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_bitslip_wait_cnt = 3'b001;
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_bitslip_wait_type = "bitslip_cnt";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_bypass = "blksync_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_clken = "blksync_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_enum_invalid_sh_cnt = "enum_invalid_sh_cnt_10g";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_knum_sh_cnt_postlock = "knum_sh_cnt_postlock_10g";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_knum_sh_cnt_prelock = "knum_sh_cnt_prelock_10g";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .blksync_pipeln = "blksync_pipeln_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .clr_errblk_cnt_en = "disable";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .control_del = "control_del_none";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .crcchk_bypass = "crcchk_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .crcchk_clken = "crcchk_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .crcchk_inv = "crcchk_inv_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .crcchk_pipeln = "crcchk_pipeln_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .crcflag_pipeln = "crcflag_pipeln_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .ctrl_bit_reverse = "ctrl_bit_reverse_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .data_bit_reverse = "data_bit_reverse_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .dec64b66b_clken = "dec64b66b_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .dec_64b66b_rxsm_bypass = "dec_64b66b_rxsm_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .descrm_bypass = "descrm_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .descrm_clken = "descrm_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .descrm_mode = "async";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .descrm_pipeln = "enable";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .dft_clk_out_sel = "rx_master_clk";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .dis_signal_ok = "dis_signal_ok_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .dispchk_bypass = "dispchk_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .empty_flag_type = "empty_rd_side";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fast_path = "fast_path_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fec_clken = "fec_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fec_enable = "fec_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fifo_double_read = "fifo_double_read_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fifo_stop_rd = "n_rd_empty";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .fifo_stop_wr = "n_wr_full";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .force_align = "force_align_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_bypass = "frmsync_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_clken = "frmsync_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_enum_scrm = "enum_scrm_default";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_enum_sync = "enum_sync_default";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_flag_type = "location_only";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_knum_sync = "knum_sync_default";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_mfrm_length = 16'b0000100000000000;
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .frmsync_pipeln = "frmsync_pipeln_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .full_flag_type = "full_wr_side";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .gb_rx_idwidth = "width_64";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .gb_rx_odwidth = "width_64";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .gbexp_clken = "gbexp_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .low_latency_en = "disable";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .lpbk_mode = "lpbk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .master_clk_sel = "master_rx_pma_clk";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .pempty_flag_type = "pempty_rd_side";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .pfull_flag_type = "pfull_wr_side";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .phcomp_rd_del = "phcomp_rd_del2";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .pld_if_type = "fifo";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .prot_mode = "disable_mode";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rand_clken = "rand_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rd_clk_sel = "rd_rx_pld_clk";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rdfifo_clken = "rdfifo_clk_dis";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_fifo_write_ctrl = "blklock_stops";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_scrm_width = "bit64";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_sh_location = "msb";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_signal_ok_sel = "synchronized_ver";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_sm_bypass = "rx_sm_bypass_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_sm_hiber = "rx_sm_hiber_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_sm_pipeln = "rx_sm_pipeln_en";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_testbus_sel = "rx_fifo_testbus1";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rx_true_b2b = "b2b";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rxfifo_empty = "empty_default";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rxfifo_full = "full_default";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rxfifo_mode = "phase_comp";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rxfifo_pempty = 5'b00010;
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .rxfifo_pfull = 5'b10111;
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .stretch_num_stages = "zero_stage";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .test_mode = "test_off";
defparam \gen_twentynm_hssi_10g_rx_pcs.inst_twentynm_hssi_10g_rx_pcs .wrfifo_clken = "wrfifo_clk_dis";

twentynm_hssi_8g_rx_pcs \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs (
	.a1a2_size(w_hssi_rx_pld_pcs_interface_int_pldif_8g_a1a2_size),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.bit_reversal_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitloc_rev_en),
	.bitslip(w_hssi_rx_pld_pcs_interface_int_pldif_8g_bitslip),
	.byte_rev_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_byte_rev_en),
	.disable_pc_fifo_byte_serdes(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[4] ),
	.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
	.eios_detected_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
	.enable_comma_detect(w_hssi_rx_pld_pcs_interface_int_pldif_8g_encdt),
	.gen3_clk_sel(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2] ),
	.hrd_rst(gnd),
	.inferred_rxvalid_cdr_ctrl(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
	.pc_fifo_rd_enable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rdenable_rx),
	.pc_fifo_wrdisable(w_hssi_rx_pld_pcs_interface_int_pldif_8g_wrdisable_rx),
	.pcie_switch(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8] ),
	.pcs_rst(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3] ),
	.phystatus_int(w_hssi_pipe_gen1_2_phystatus),
	.phystatus_pcs_gen3(w_hssi_pipe_gen3_phystatus),
	.pipe_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
	.pld_rx_clk(w_hssi_rx_pld_pcs_interface_int_pldif_8g_pld_rx_clk),
	.polarity_inversion(w_hssi_pipe_gen1_2_polarity_inversion_rx),
	.rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
	.rd_enable_in_chnl_down(gnd),
	.rd_enable_in_chnl_up(gnd),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
	.refclk_dig2(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig2),
	.reset_pc_ptrs_asn(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[5] ),
	.reset_pc_ptrs_in_chnl_down(gnd),
	.reset_pc_ptrs_in_chnl_up(gnd),
	.reset_ppm_cntrs_pcs_pma(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[7] ),
	.rm_fifo_read_enable(gnd),
	.rm_fifo_write_enable(gnd),
	.rx_pcs_rst(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxurstpcs_n),
	.rxvalid_int(w_hssi_pipe_gen1_2_rxvalid),
	.rxvalid_pcs_gen3(w_hssi_pipe_gen3_rxvalid),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
	.sig_det_from_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
	.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
	.speed_change(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0] ),
	.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
	.syncsm_en(w_hssi_rx_pld_pcs_interface_int_pldif_8g_syncsm_en),
	.tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
	.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
	.wr_enable_in_chnl_down(gnd),
	.wr_enable_in_chnl_up(gnd),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.datain({\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[19] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[18] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[17] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[16] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[15] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[14] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[13] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[12] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[11] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[10] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[9] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[8] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[7] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[6] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[5] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[4] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[3] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[2] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[1] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_8g_pudi[0] }),
	.eidleinfersel({\w_hssi_8g_tx_pcs_non_gray_eidleinfersel[2] ,\w_hssi_8g_tx_pcs_non_gray_eidleinfersel[1] ,\w_hssi_8g_tx_pcs_non_gray_eidleinfersel[0] }),
	.rd_data1_rx_rmfifo({\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[31] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[30] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[29] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[28] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[27] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[26] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[25] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[24] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[23] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[22] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[21] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[20] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[19] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[18] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[17] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[16] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[15] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[14] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[13] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[12] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[11] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[10] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[9] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[8] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[7] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[6] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[5] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[4] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[3] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[2] ,
\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[1] ,\w_hssi_fifo_rx_pcs_data_out_8g_clock_comp[0] }),
	.rd_data2_rx_rmfifo({\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[31] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[30] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[29] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[28] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[27] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[26] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[25] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[24] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[23] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[22] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[21] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[20] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[19] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[18] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[17] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[16] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[15] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[14] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[13] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[12] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[11] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[10] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[9] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[8] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[7] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[6] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[5] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[4] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[3] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[2] ,
\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[1] ,\w_hssi_fifo_rx_pcs_data_out2_8g_clock_comp[0] }),
	.rd_data_rx_phfifo({\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[79] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[78] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[77] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[76] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[75] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[74] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[73] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[72] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[71] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[70] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[69] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[68] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[67] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[66] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[65] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[64] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[63] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[62] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[61] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[60] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[59] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[58] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[57] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[56] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[55] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[54] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[53] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[52] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[51] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[50] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[49] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[48] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[47] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[46] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[45] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[44] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[43] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[42] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[41] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[40] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[39] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[38] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[37] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[36] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[35] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[34] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[33] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[32] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[31] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[30] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[29] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[28] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[27] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[26] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[25] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[24] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[23] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[22] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[21] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[20] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[19] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[18] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[17] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[16] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[15] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[14] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[13] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[12] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[11] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[10] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[9] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[8] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[7] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[6] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[5] ,
\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[4] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[3] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[2] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[1] ,\w_hssi_fifo_rx_pcs_data_out_8g_phase_comp[0] }),
	.rx_blk_start_pcs_gen3({\w_hssi_pipe_gen3_rx_blk_start[3] ,\w_hssi_pipe_gen3_rx_blk_start[2] ,\w_hssi_pipe_gen3_rx_blk_start[1] ,\w_hssi_pipe_gen3_rx_blk_start[0] }),
	.rx_data_pcs_gen3({\w_hssi_pipe_gen3_rxd_8gpcs_out[63] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[62] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[61] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[60] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[59] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[58] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[57] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[56] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[55] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[54] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[53] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[52] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[51] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[50] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[49] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[48] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[47] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[46] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[45] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[44] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[43] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[42] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[41] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[40] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[39] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[38] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[37] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[36] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[35] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[34] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[33] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[32] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[31] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[30] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[29] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[28] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[27] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[26] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[25] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[24] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[23] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[22] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[21] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[20] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[19] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[18] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[17] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[16] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[15] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[14] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[13] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[12] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[11] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[10] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[9] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[8] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[7] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[6] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[5] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[4] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[3] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[2] ,\w_hssi_pipe_gen3_rxd_8gpcs_out[1] ,
\w_hssi_pipe_gen3_rxd_8gpcs_out[0] }),
	.rx_data_valid_pcs_gen3({\w_hssi_pipe_gen3_rxdataskip[3] ,\w_hssi_pipe_gen3_rxdataskip[2] ,\w_hssi_pipe_gen3_rxdataskip[1] ,\w_hssi_pipe_gen3_rxdataskip[0] }),
	.rx_div_sync_in_chnl_down({gnd,gnd}),
	.rx_div_sync_in_chnl_up({gnd,gnd}),
	.rx_sync_hdr_pcs_gen3({\w_hssi_pipe_gen3_rx_sync_hdr[1] ,\w_hssi_pipe_gen3_rx_sync_hdr[0] }),
	.rx_we_in_chnl_down({gnd,gnd}),
	.rx_we_in_chnl_up({gnd,gnd}),
	.rxstatus_int({\w_hssi_pipe_gen1_2_rxstatus[2] ,\w_hssi_pipe_gen1_2_rxstatus[1] ,\w_hssi_pipe_gen1_2_rxstatus[0] }),
	.rxstatus_pcs_gen3({\w_hssi_pipe_gen3_rxstatus[2] ,\w_hssi_pipe_gen3_rxstatus[1] ,\w_hssi_pipe_gen3_rxstatus[0] }),
	.tx_ctrlplane_testbus({\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[19] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[18] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[17] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[16] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[15] ,
\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[14] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[13] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[12] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[11] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[10] ,
\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[9] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[8] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[7] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[6] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[5] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[4] ,
\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[3] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[2] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[1] ,\w_hssi_8g_tx_pcs_tx_ctrlplane_testbus[0] }),
	.tx_div_sync({\w_hssi_8g_tx_pcs_tx_div_sync[1] ,\w_hssi_8g_tx_pcs_tx_div_sync[0] }),
	.tx_testbus({\w_hssi_8g_tx_pcs_tx_testbus[19] ,\w_hssi_8g_tx_pcs_tx_testbus[18] ,\w_hssi_8g_tx_pcs_tx_testbus[17] ,\w_hssi_8g_tx_pcs_tx_testbus[16] ,\w_hssi_8g_tx_pcs_tx_testbus[15] ,\w_hssi_8g_tx_pcs_tx_testbus[14] ,\w_hssi_8g_tx_pcs_tx_testbus[13] ,
\w_hssi_8g_tx_pcs_tx_testbus[12] ,\w_hssi_8g_tx_pcs_tx_testbus[11] ,\w_hssi_8g_tx_pcs_tx_testbus[10] ,\w_hssi_8g_tx_pcs_tx_testbus[9] ,\w_hssi_8g_tx_pcs_tx_testbus[8] ,\w_hssi_8g_tx_pcs_tx_testbus[7] ,\w_hssi_8g_tx_pcs_tx_testbus[6] ,
\w_hssi_8g_tx_pcs_tx_testbus[5] ,\w_hssi_8g_tx_pcs_tx_testbus[4] ,\w_hssi_8g_tx_pcs_tx_testbus[3] ,\w_hssi_8g_tx_pcs_tx_testbus[2] ,\w_hssi_8g_tx_pcs_tx_testbus[1] ,\w_hssi_8g_tx_pcs_tx_testbus[0] }),
	.blockselect(out_blockselect_hssi_8g_rx_pcs),
	.byte_deserializer_pcs_clk_div_by_2_reg(),
	.byte_deserializer_pcs_clk_div_by_2_txclk_reg(),
	.byte_deserializer_pcs_clk_div_by_2_txclk_wire(),
	.byte_deserializer_pcs_clk_div_by_2_wire(),
	.byte_deserializer_pcs_clk_div_by_4_txclk_reg(),
	.byte_deserializer_pld_clk_div_by_2_reg(),
	.byte_deserializer_pld_clk_div_by_2_txclk_reg(),
	.byte_deserializer_pld_clk_div_by_4_txclk_reg(),
	.clock_to_pld(w_hssi_8g_rx_pcs_clock_to_pld),
	.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
	.eidle_detected(w_hssi_8g_rx_pcs_eidle_detected),
	.g3_rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
	.g3_rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
	.gen2ngen1(w_hssi_8g_rx_pcs_gen2ngen1),
	.pc_fifo_empty(w_hssi_8g_rx_pcs_pc_fifo_empty),
	.pcfifofull(w_hssi_8g_rx_pcs_pcfifofull),
	.phystatus(w_hssi_8g_rx_pcs_phystatus),
	.pld_8g_a1a2_k1k2_flag_reg(),
	.pld_8g_a1a2_k1k2_flag_txclk_reg(),
	.pld_8g_a1a2_size_reg(),
	.pld_8g_a1a2_size_txclk_reg(),
	.pld_8g_bitloc_rev_en_reg(),
	.pld_8g_bitloc_rev_en_txclk_reg(),
	.pld_8g_byte_rev_en_reg(),
	.pld_8g_byte_rev_en_txclk_reg(),
	.pld_8g_elecidle_reg(),
	.pld_8g_empty_rmf_lowlatency_reg(),
	.pld_8g_empty_rmf_lowlatency_txclk_reg(),
	.pld_8g_empty_rmf_reg(),
	.pld_8g_empty_rmf_txclk_reg(),
	.pld_8g_empty_rx_fifo(),
	.pld_8g_empty_rx_reg(),
	.pld_8g_empty_rx_txclk_reg(),
	.pld_8g_encdt_reg(),
	.pld_8g_encdt_txclk_reg(),
	.pld_8g_full_rmf_reg(),
	.pld_8g_full_rmf_txclk_reg(),
	.pld_8g_full_rx_fifo(),
	.pld_8g_full_rx_reg(),
	.pld_8g_full_rx_txclk_reg(),
	.pld_8g_g3_rx_pld_rst_n_reg(),
	.pld_8g_g3_rx_pld_rst_n_txclk_reg(),
	.pld_8g_rxelecidle_txclk_reg(),
	.pld_8g_rxpolarity_reg(),
	.pld_8g_rxpolarity_txclk_reg(),
	.pld_8g_wa_boundary_reg(),
	.pld_8g_wrdisable_rx_reg(),
	.pld_8g_wrdisable_rx_txclk_reg(),
	.pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire(),
	.pld_pcs_rx_clk_out_8g_div_by_2_wire(),
	.pld_pcs_rx_clk_out_8g_txclk_wire(),
	.pld_pcs_rx_clk_out_8g_wire(),
	.pld_rx_control_8g_reg(),
	.pld_rx_control_8g_txclk_reg(),
	.pld_rx_data_8g_reg(),
	.pld_rx_data_8g_txclk_reg(),
	.pld_syncsm_en_reg(),
	.pld_syncsm_en_txclk_reg(),
	.rd_enable_out_chnl_down(),
	.rd_enable_out_chnl_up(),
	.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
	.reset_pc_ptrs_in_chnl_down_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
	.reset_pc_ptrs_in_chnl_up_pipe(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
	.reset_pc_ptrs_out_chnl_down(),
	.reset_pc_ptrs_out_chnl_up(),
	.rm_fifo_empty(w_hssi_8g_rx_pcs_rm_fifo_empty),
	.rm_fifo_full(w_hssi_8g_rx_pcs_rm_fifo_full),
	.rm_fifo_partial_empty(),
	.rm_fifo_partial_full(),
	.rx_clk_out_pld_if(w_hssi_8g_rx_pcs_rx_clk_out_pld_if),
	.rx_clk_to_observation_ff_in_pld_if(w_hssi_8g_rx_pcs_rx_clk_to_observation_ff_in_pld_if),
	.rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
	.rx_pipe_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
	.rx_pipe_soft_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
	.rx_pma_clk_gen3(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
	.rx_rcvd_clk_gen3(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
	.rx_rstn_sync2wrfifo_8g(w_hssi_8g_rx_pcs_rx_rstn_sync2wrfifo_8g),
	.rxvalid(w_hssi_8g_rx_pcs_rxvalid),
	.signal_detect_out(w_hssi_8g_rx_pcs_signal_detect_out),
	.sta_rx_clk2_by2_1(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs~O_STA_RX_CLK2_BY2_1 ),
	.sta_rx_clk2_by2_1_out(),
	.sta_rx_clk2_by2_2(),
	.sta_rx_clk2_by2_2_out(),
	.sta_rx_clk2_by4_1(),
	.sta_rx_clk2_by4_1_out(),
	.wr_clk_rx_phfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
	.wr_clk_rx_phfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
	.wr_clk_rx_rmfifo_dw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
	.wr_clk_rx_rmfifo_sw_clk(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
	.wr_en_rx_phfifo(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
	.wr_en_rx_rmfifo(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
	.wr_enable_out_chnl_down(),
	.wr_enable_out_chnl_up(),
	.wr_rst_n_rx_phfifo(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
	.wr_rst_rx_rmfifo(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
	.a1a2k1k2flag(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_A1A2K1K2FLAG_bus ),
	.avmmreaddata(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_AVMMREADDATA_bus ),
	.chnl_test_bus_out(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_CHNL_TEST_BUS_OUT_bus ),
	.dataout(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_DATAOUT_bus ),
	.eios_det_cdr_ctrl(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_EIOS_DET_CDR_CTRL_bus ),
	.parallel_rev_loopback(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PARALLEL_REV_LOOPBACK_bus ),
	.pipe_data(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_PIPE_DATA_bus ),
	.rd_ptr1_rx_rmfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR1_RX_RMFIFO_bus ),
	.rd_ptr2_rx_rmfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR2_RX_RMFIFO_bus ),
	.rd_ptr_rx_phfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RD_PTR_RX_PHFIFO_bus ),
	.rx_blk_start(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_BLK_START_bus ),
	.rx_data_valid(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_DATA_VALID_bus ),
	.rx_div_sync_out_chnl_down(),
	.rx_div_sync_out_chnl_up(),
	.rx_sync_hdr(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RX_SYNC_HDR_bus ),
	.rx_we_out_chnl_down(),
	.rx_we_out_chnl_up(),
	.rxstatus(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_RXSTATUS_bus ),
	.word_align_boundary(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WORD_ALIGN_BOUNDARY_bus ),
	.wr_data_rx_phfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_PHFIFO_bus ),
	.wr_data_rx_rmfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_DATA_RX_RMFIFO_bus ),
	.wr_ptr_rx_phfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_PHFIFO_bus ),
	.wr_ptr_rx_rmfifo(\gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs_WR_PTR_RX_RMFIFO_bus ));
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .auto_error_replacement = "dis_err_replace";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .auto_speed_nego = "dis_asn";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .bit_reversal = "dis_bit_reversal";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .bonding_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .bonding_dft_val = "dft_0";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .bypass_pipeline_reg = "dis_bypass_pipeline";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .byte_deserializer = "dis_bds";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .cdr_ctrl_rxvalid_mask = "dis_rxvalid_mask";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clkcmp_pattern_n = 20'b00000000000000000000;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clkcmp_pattern_p = 20'b00000000000000000000;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_bds_dec_asn = "dis_bds_dec_asn_clk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_cdr_eidle = "en_cdr_eidle_clk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_dw_pc_wrclk = "en_dw_pc_wrclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_dw_rm_rd = "en_dw_rm_rdclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_dw_rm_wr = "en_dw_rm_wrclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_dw_wa = "en_dw_wa_clk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_pc_rdclk = "dis_pc_rdclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_sw_pc_wrclk = "dis_sw_pc_wrclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_sw_rm_rd = "en_sw_rm_rdclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_sw_rm_wr = "en_sw_rm_wrclk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_gate_sw_wa = "dis_sw_wa_clk_gating";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .clock_observation_in_pld_core = "internal_sw_wa_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .ctrl_plane_bonding_compensation = "dis_compensation";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .ctrl_plane_bonding_consumption = "individual";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .ctrl_plane_bonding_distribution = "not_master_chnl_distr";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .eidle_entry_eios = "dis_eidle_eios";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .eidle_entry_iei = "dis_eidle_iei";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .eidle_entry_sd = "dis_eidle_sd";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .eightb_tenb_decoder = "en_8b10b_ibm";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .err_flags_sel = "err_flags_wa";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .fixed_pat_det = "dis_fixed_patdet";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .fixed_pat_num = 4'b0000;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .force_signal_detect = "en_force_signal_detect";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .gen3_clk_en = "disable_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .gen3_rx_clk_sel = "rcvd_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .gen3_tx_clk_sel = "tx_pma_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .hip_mode = "dis_hip";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .ibm_invalid_code = "dis_ibm_invalid_code";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .invalid_code_flag_only = "dis_invalid_code_only";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .pad_or_edb_error_replace = "replace_edb";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .pcs_bypass = "dis_pcs_bypass";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .phase_comp_rdptr = "disable_rdptr";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .phase_compensation_fifo = "register_fifo";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .pipe_if_enable = "dis_pipe_rx";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .pma_dw = "ten_bit";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .polinv_8b10b_dec = "dis_polinv_8b10b_dec";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .prot_mode = "cpri_rx_tx";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match = "dis_rm";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match_del_thres = "dis_rm_del_thres";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match_empty_thres = "dis_rm_empty_thres";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match_full_thres = "dis_rm_full_thres";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match_ins_thres = "dis_rm_ins_thres";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rate_match_start_thres = "dis_rm_start_thres";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_clk2 = "rcvd_clk_clk2";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_clk_free_running = "en_rx_clk_free_run";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_pcs_urst = "en_rx_pcs_urst";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_rcvd_clk = "rcvd_clk_rcvd_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_rd_clk = "rx_clk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_refclk = "dis_refclk_sel";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .rx_wr_clk = "rx_clk2_div_1_2_4";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .symbol_swap = "dis_symbol_swap";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .sync_sm_idle_eios = "dis_syncsm_idle";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .test_bus_sel = "tx_testbus";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .tx_rx_parallel_loopback = "dis_plpbk";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_boundary_lock_ctrl = "auto_align_pld_ctrl";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_clk_slip_spacing = 10'b0000010000;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_det_latency_sync_status_beh = "dont_care_assert_sync";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_disp_err_flag = "en_disp_err_flag";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_kchar = "dis_kchar";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_pd = "wa_pd_10";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_pd_data = 40'b0000000000000000000000000000000101111100;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_pd_polarity = "dont_care_both_pol";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_pld_controlled = "pld_ctrl_sw";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_renumber_data = 6'b000011;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_rgnumber_data = 8'b00000011;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_rknumber_data = 8'b00000011;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_rosnumber_data = 2'b01;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_rvnumber_data = 13'b0000000000000;
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wa_sync_sm_ctrl = "gige_sync_sm";
defparam \gen_twentynm_hssi_8g_rx_pcs.inst_twentynm_hssi_8g_rx_pcs .wait_cnt = 12'b000000000000;

twentynm_hssi_pipe_gen1_2 \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.pcie_switch(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[8] ),
	.pipe_rx_clk(w_hssi_8g_rx_pcs_rx_pipe_clk),
	.pipe_tx_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
	.power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
	.power_state_transition_done_ena(gnd),
	.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
	.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
	.rev_loopbk_pcs_gen3(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
	.revloopback(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
	.rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
	.rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
	.rx_pipe_reset(w_hssi_8g_rx_pcs_rx_pipe_soft_reset),
	.rxelectricalidle(w_hssi_8g_rx_pcs_eidle_detected),
	.rxelectricalidle_pcs_gen3(w_hssi_pipe_gen3_rxelecidle),
	.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
	.rxpolarity_pcs_gen3(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
	.sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
	.speed_change(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[0] ),
	.tx_elec_idle_comp(w_hssi_8g_tx_pcs_tx_pipe_electidle),
	.tx_pipe_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
	.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
	.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
	.txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txelecidle),
	.txswingport(w_hssi_8g_tx_pcs_phfifo_txswing),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.powerdown({\w_hssi_8g_tx_pcs_pipe_power_down_out[1] ,\w_hssi_8g_tx_pcs_pipe_power_down_out[0] }),
	.rxd({\w_hssi_8g_rx_pcs_pipe_data[63] ,\w_hssi_8g_rx_pcs_pipe_data[62] ,\w_hssi_8g_rx_pcs_pipe_data[61] ,\w_hssi_8g_rx_pcs_pipe_data[60] ,\w_hssi_8g_rx_pcs_pipe_data[59] ,\w_hssi_8g_rx_pcs_pipe_data[58] ,\w_hssi_8g_rx_pcs_pipe_data[57] ,\w_hssi_8g_rx_pcs_pipe_data[56] ,
\w_hssi_8g_rx_pcs_pipe_data[55] ,\w_hssi_8g_rx_pcs_pipe_data[54] ,\w_hssi_8g_rx_pcs_pipe_data[53] ,\w_hssi_8g_rx_pcs_pipe_data[52] ,\w_hssi_8g_rx_pcs_pipe_data[51] ,\w_hssi_8g_rx_pcs_pipe_data[50] ,\w_hssi_8g_rx_pcs_pipe_data[49] ,\w_hssi_8g_rx_pcs_pipe_data[48] ,
\w_hssi_8g_rx_pcs_pipe_data[47] ,\w_hssi_8g_rx_pcs_pipe_data[46] ,\w_hssi_8g_rx_pcs_pipe_data[45] ,\w_hssi_8g_rx_pcs_pipe_data[44] ,\w_hssi_8g_rx_pcs_pipe_data[43] ,\w_hssi_8g_rx_pcs_pipe_data[42] ,\w_hssi_8g_rx_pcs_pipe_data[41] ,\w_hssi_8g_rx_pcs_pipe_data[40] ,
\w_hssi_8g_rx_pcs_pipe_data[39] ,\w_hssi_8g_rx_pcs_pipe_data[38] ,\w_hssi_8g_rx_pcs_pipe_data[37] ,\w_hssi_8g_rx_pcs_pipe_data[36] ,\w_hssi_8g_rx_pcs_pipe_data[35] ,\w_hssi_8g_rx_pcs_pipe_data[34] ,\w_hssi_8g_rx_pcs_pipe_data[33] ,\w_hssi_8g_rx_pcs_pipe_data[32] ,
\w_hssi_8g_rx_pcs_pipe_data[31] ,\w_hssi_8g_rx_pcs_pipe_data[30] ,\w_hssi_8g_rx_pcs_pipe_data[29] ,\w_hssi_8g_rx_pcs_pipe_data[28] ,\w_hssi_8g_rx_pcs_pipe_data[27] ,\w_hssi_8g_rx_pcs_pipe_data[26] ,\w_hssi_8g_rx_pcs_pipe_data[25] ,\w_hssi_8g_rx_pcs_pipe_data[24] ,
\w_hssi_8g_rx_pcs_pipe_data[23] ,\w_hssi_8g_rx_pcs_pipe_data[22] ,\w_hssi_8g_rx_pcs_pipe_data[21] ,\w_hssi_8g_rx_pcs_pipe_data[20] ,\w_hssi_8g_rx_pcs_pipe_data[19] ,\w_hssi_8g_rx_pcs_pipe_data[18] ,\w_hssi_8g_rx_pcs_pipe_data[17] ,\w_hssi_8g_rx_pcs_pipe_data[16] ,
\w_hssi_8g_rx_pcs_pipe_data[15] ,\w_hssi_8g_rx_pcs_pipe_data[14] ,\w_hssi_8g_rx_pcs_pipe_data[13] ,\w_hssi_8g_rx_pcs_pipe_data[12] ,\w_hssi_8g_rx_pcs_pipe_data[11] ,\w_hssi_8g_rx_pcs_pipe_data[10] ,\w_hssi_8g_rx_pcs_pipe_data[9] ,\w_hssi_8g_rx_pcs_pipe_data[8] ,
\w_hssi_8g_rx_pcs_pipe_data[7] ,\w_hssi_8g_rx_pcs_pipe_data[6] ,\w_hssi_8g_rx_pcs_pipe_data[5] ,\w_hssi_8g_rx_pcs_pipe_data[4] ,\w_hssi_8g_rx_pcs_pipe_data[3] ,\w_hssi_8g_rx_pcs_pipe_data[2] ,\w_hssi_8g_rx_pcs_pipe_data[1] ,\w_hssi_8g_rx_pcs_pipe_data[0] }),
	.txd_ch({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0] }),
	.txmargin({\w_hssi_8g_tx_pcs_phfifo_txmargin[2] ,\w_hssi_8g_tx_pcs_phfifo_txmargin[1] ,\w_hssi_8g_tx_pcs_phfifo_txmargin[0] }),
	.blockselect(out_blockselect_hssi_pipe_gen1_2),
	.phystatus(w_hssi_pipe_gen1_2_phystatus),
	.pld_8g_rxpolarity_pipe3_reg(),
	.polarity_inversion_rx(w_hssi_pipe_gen1_2_polarity_inversion_rx),
	.rev_loopbk(w_hssi_pipe_gen1_2_rev_loopbk),
	.rxelecidle(w_hssi_pipe_gen1_2_rxelecidle),
	.rxelectricalidle_out(w_hssi_pipe_gen1_2_rxelectricalidle_out),
	.rxvalid(w_hssi_pipe_gen1_2_rxvalid),
	.tx_elec_idle_out(w_hssi_pipe_gen1_2_tx_elec_idle_out),
	.txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
	.avmmreaddata(\gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_AVMMREADDATA_bus ),
	.current_coeff(\gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_CURRENT_COEFF_bus ),
	.rxd_ch(),
	.rxstatus(\gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2_RXSTATUS_bus ),
	.txd());
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .elec_idle_delay_val = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .error_replace_pad = "replace_edb";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .hip_mode = "dis_hip";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .ind_error_reporting = "dis_ind_error_reporting";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .phystatus_delay_val = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .phystatus_rst_toggle = "dis_phystatus_rst_toggle";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .pipe_byte_de_serializer_en = "dont_care_bds";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .prot_mode = "disabled_prot_mode";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rpre_emph_a_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rpre_emph_b_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rpre_emph_c_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rpre_emph_d_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rpre_emph_e_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rvod_sel_a_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rvod_sel_b_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rvod_sel_c_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rvod_sel_d_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rvod_sel_e_val = 6'b000000;
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rx_pipe_enable = "dis_pipe_rx";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .rxdetect_bypass = "dis_rxdetect_bypass";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .tx_pipe_enable = "dis_pipe_tx";
defparam \gen_twentynm_hssi_pipe_gen1_2.inst_twentynm_hssi_pipe_gen1_2 .txswing = "dis_txswing";

twentynm_hssi_krfec_rx_pcs \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.rx_clr_counters(w_hssi_rx_pld_pcs_interface_int_pldif_krfec_rx_clr_counters),
	.rx_krfec_clk(w_hssi_10g_rx_pcs_rx_fec_clk),
	.rx_master_clk(w_hssi_10g_rx_pcs_rx_master_clk),
	.rx_master_clk_rst_n(w_hssi_10g_rx_pcs_rx_master_clk_rst_n),
	.rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_mode_n),
	.scan_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_krfec_scan_rst_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.rx_data_in({\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[63] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[62] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[61] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[60] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[59] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[58] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[57] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[56] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[55] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[54] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[53] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[52] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[51] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[50] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[49] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[48] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[47] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[46] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[45] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[44] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[43] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[42] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[41] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[40] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[39] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[38] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[37] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[36] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[35] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[34] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[33] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[32] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[31] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[30] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[29] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[28] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[27] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[26] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[25] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[24] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[23] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[22] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[21] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[20] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[19] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[18] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[17] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[16] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[15] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[14] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[13] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[12] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[11] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[10] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[9] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[8] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[7] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[6] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[5] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[4] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[3] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[2] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[1] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_pma_data[0] }),
	.blockselect(out_blockselect_hssi_krfec_rx_pcs),
	.pld_10g_krfec_rx_blk_lock_krfec_reg(),
	.pld_10g_krfec_rx_blk_lock_krfec_txclk_reg(),
	.pld_10g_krfec_rx_diag_data_status_krfec_reg(),
	.pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg(),
	.pld_10g_krfec_rx_frame_krfec_reg(),
	.pld_10g_krfec_rx_frame_krfec_txclk_reg(),
	.rx_block_lock(w_hssi_krfec_rx_pcs_rx_block_lock),
	.rx_data_valid_out(w_hssi_krfec_rx_pcs_rx_data_valid_out),
	.rx_frame(w_hssi_krfec_rx_pcs_rx_frame),
	.rx_signal_ok_out(w_hssi_krfec_rx_pcs_rx_signal_ok_out),
	.avmmreaddata(\gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_AVMMREADDATA_bus ),
	.rx_control_out(\gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_CONTROL_OUT_bus ),
	.rx_data_out(\gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_OUT_bus ),
	.rx_data_status(\gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs_RX_DATA_STATUS_bus ),
	.rx_test_data());
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .blksync_cor_en = "detect";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .bypass_gb = "bypass_dis";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .clr_ctrl = "both_enabled";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .ctrl_bit_reverse = "ctrl_bit_reverse_en";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .data_bit_reverse = "data_bit_reverse_dis";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .dv_start = "with_blklock";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .err_mark_type = "err_mark_10g";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .error_marking_en = "err_mark_dis";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .low_latency_en = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .lpbk_mode = "lpbk_dis";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .parity_invalid_enum = 8'b00001000;
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .parity_valid_num = 4'b0100;
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_blksync = "enable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_descrm = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_errcorrect = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_errtrap_ind = "enable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_errtrap_lfsr = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_errtrap_loc = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_errtrap_pat = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_gearbox = "enable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_syndrm = "enable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .pipeln_trans_dec = "disable";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .prot_mode = "disable_mode";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .receive_order = "receive_lsb";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .rx_testbus_sel = "overall";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .signal_ok_en = "sig_ok_en";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_krfec_rx_pcs.inst_twentynm_hssi_krfec_rx_pcs .sup_mode = "user_mode";

twentynm_hssi_rx_pcs_pma_interface \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pmaif_10g_random_err(w_hssi_10g_rx_pcs_rx_random_err),
	.int_pmaif_8g_rx_clkslip(w_hssi_8g_rx_pcs_rx_clkslip),
	.int_pmaif_pldif_pmaif_rx_pld_rst_n(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_pld_rst_n),
	.int_pmaif_pldif_polinv_rx(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_polinv_rx),
	.int_pmaif_pldif_prbs_err_clr(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_prbs_err_clr),
	.int_pmaif_pldif_rx_clkslip(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rx_clkslip),
	.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
	.pma_rx_clkdiv_user(in_pma_rx_clkdiv_user),
	.pma_rx_detect_valid(in_pma_rx_detect_valid),
	.pma_rx_found(in_pma_rx_found),
	.pma_rx_pma_clk(in_pma_rx_pma_clk),
	.pma_rx_signal_ok(vcc),
	.pma_rxpll_lock(in_pma_rxpll_lock),
	.pma_signal_det(in_pma_signal_det),
	.pma_tx_pma_clk(in_pma_tx_pma_clk),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.int_pmaif_pldif_eye_monitor({\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[5] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[4] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[3] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[2] ,
\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_eye_monitor[0] }),
	.pma_rx_pma_data({in_pma_rx_pma_data[63],in_pma_rx_pma_data[62],in_pma_rx_pma_data[61],in_pma_rx_pma_data[60],in_pma_rx_pma_data[59],in_pma_rx_pma_data[58],in_pma_rx_pma_data[57],in_pma_rx_pma_data[56],in_pma_rx_pma_data[55],in_pma_rx_pma_data[54],in_pma_rx_pma_data[53],in_pma_rx_pma_data[52],in_pma_rx_pma_data[51],in_pma_rx_pma_data[50],
in_pma_rx_pma_data[49],in_pma_rx_pma_data[48],in_pma_rx_pma_data[47],in_pma_rx_pma_data[46],in_pma_rx_pma_data[45],in_pma_rx_pma_data[44],in_pma_rx_pma_data[43],in_pma_rx_pma_data[42],in_pma_rx_pma_data[41],in_pma_rx_pma_data[40],in_pma_rx_pma_data[39],in_pma_rx_pma_data[38],in_pma_rx_pma_data[37],in_pma_rx_pma_data[36],
in_pma_rx_pma_data[35],in_pma_rx_pma_data[34],in_pma_rx_pma_data[33],in_pma_rx_pma_data[32],in_pma_rx_pma_data[31],in_pma_rx_pma_data[30],in_pma_rx_pma_data[29],in_pma_rx_pma_data[28],in_pma_rx_pma_data[27],in_pma_rx_pma_data[26],in_pma_rx_pma_data[25],in_pma_rx_pma_data[24],in_pma_rx_pma_data[23],in_pma_rx_pma_data[22],
in_pma_rx_pma_data[21],in_pma_rx_pma_data[20],in_pma_rx_pma_data[19],in_pma_rx_pma_data[18],in_pma_rx_pma_data[17],in_pma_rx_pma_data[16],in_pma_rx_pma_data[15],in_pma_rx_pma_data[14],in_pma_rx_pma_data[13],in_pma_rx_pma_data[12],in_pma_rx_pma_data[11],in_pma_rx_pma_data[10],in_pma_rx_pma_data[9],in_pma_rx_pma_data[8],
in_pma_rx_pma_data[7],in_pma_rx_pma_data[6],in_pma_rx_pma_data[5],in_pma_rx_pma_data[4],in_pma_rx_pma_data[3],in_pma_rx_pma_data[2],in_pma_rx_pma_data[1],in_pma_rx_pma_data[0]}),
	.tx_pma_data_loopback({\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[63] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[62] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[61] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[60] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[59] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[58] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[57] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[56] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[55] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[54] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[53] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[52] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[51] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[50] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[49] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[48] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[47] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[46] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[45] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[44] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[43] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[42] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[41] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[40] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[39] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[38] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[37] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[36] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[35] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[34] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[33] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[32] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[31] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[30] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[29] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[28] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[27] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[26] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[25] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[24] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[23] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[22] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[21] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[20] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[19] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[18] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[17] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[16] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[15] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[14] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[13] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[12] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[11] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[10] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[9] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[8] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[7] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[6] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[5] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[4] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[3] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[2] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[1] ,\w_hssi_tx_pcs_pma_interface_tx_pma_data_loopback[0] }),
	.tx_pma_uhsif_data_loopback({\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[63] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[62] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[61] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[60] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[59] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[58] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[57] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[56] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[55] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[54] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[53] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[52] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[51] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[50] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[49] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[48] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[47] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[46] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[45] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[44] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[43] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[42] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[41] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[40] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[39] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[38] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[37] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[36] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[35] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[34] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[33] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[32] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[31] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[30] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[29] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[28] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[27] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[26] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[25] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[24] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[23] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[22] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[21] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[20] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[19] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[18] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[17] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[16] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[15] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[14] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[13] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[12] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[11] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[10] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[9] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[8] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[7] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[6] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[5] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[4] ,
\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[3] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[2] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[1] ,\w_hssi_tx_pcs_pma_interface_tx_pma_uhsif_data_loopback[0] }),
	.blockselect(out_blockselect_hssi_rx_pcs_pma_interface),
	.int_pmaif_10g_rx_pma_clk(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_rx_pma_clk),
	.int_pmaif_10g_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_10g_signal_ok),
	.int_pmaif_8g_rcvd_clk_pma(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rcvd_clk_pma),
	.int_pmaif_8g_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_detect_valid),
	.int_pmaif_8g_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_rx_found),
	.int_pmaif_8g_sigdetni(w_hssi_rx_pcs_pma_interface_int_pmaif_8g_sigdetni),
	.int_pmaif_g3_pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
	.int_pmaif_g3_pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
	.int_pmaif_g3_pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
	.int_pmaif_g3_rcvd_clk(),
	.int_pmaif_krfec_rx_signal_ok_in(w_hssi_rx_pcs_pma_interface_int_pmaif_krfec_rx_signal_ok_in),
	.int_pmaif_pldif_prbs_err(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err),
	.int_pmaif_pldif_prbs_err_done(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_prbs_err_done),
	.int_pmaif_pldif_rx_clkdiv(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv),
	.int_pmaif_pldif_rx_clkdiv_user(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_clkdiv_user),
	.int_pmaif_pldif_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_detect_valid),
	.int_pmaif_pldif_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rx_found),
	.int_pmaif_pldif_rxpll_lock(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_rxpll_lock),
	.int_pmaif_pldif_signal_ok(w_hssi_rx_pcs_pma_interface_int_pmaif_pldif_signal_ok),
	.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
	.pma_rx_clkslip(out_pma_rx_clkslip),
	.pma_rxpma_rstb(out_pma_rxpma_rstb),
	.prbs_err_lt(),
	.avmmreaddata(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_AVMMREADDATA_bus ),
	.int_pmaif_10g_rx_pma_data(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_10G_RX_PMA_DATA_bus ),
	.int_pmaif_8g_pudi(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_8G_PUDI_bus ),
	.int_pmaif_g3_pma_data_in(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_G3_PMA_DATA_IN_bus ),
	.int_pmaif_krfec_rx_pma_data(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_KRFEC_RX_PMA_DATA_bus ),
	.int_pmaif_pldif_rx_data(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_INT_PMAIF_PLDIF_RX_DATA_bus ),
	.pma_eye_monitor(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_PMA_EYE_MONITOR_bus ),
	.rx_pmaif_test_out(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PMAIF_TEST_OUT_bus ),
	.rx_prbs_ver_test(\gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface_RX_PRBS_VER_TEST_bus ));
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .block_sel = "eight_g_pcs";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .clkslip_sel = "pld";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .lpbk_en = "disable";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .master_clk_sel = "master_rx_pma_clk";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .pldif_datawidth_mode = "pldif_data_10bit";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .pma_dw_rx = "pma_10b_rx";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .pma_if_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .pma_if_dft_val = "dft_0";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .prbs9_dwidth = "prbs9_64b";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .prbs_clken = "prbs_clk_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .prbs_ver = "prbs_off";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .prot_mode_rx = "eightg_only_pld_mode_rx";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_dyn_polarity_inversion = "rx_dyn_polinv_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_lpbk_en = "lpbk_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_prbs_force_signal_ok = "force_sig_ok";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_prbs_mask = "prbsmask128";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_prbs_mode = "teng_mode";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_signalok_signaldet_sel = "sel_sig_det";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_static_polarity_inversion = "rx_stat_polinv_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .rx_uhsif_lpbk_en = "uhsif_lpbk_dis";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_rx_pcs_pma_interface.inst_twentynm_hssi_rx_pcs_pma_interface .sup_mode = "user_mode";

twentynm_hssi_8g_tx_pcs \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk_sel_gen3(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[2] ),
	.coreclk(w_hssi_tx_pld_pcs_interface_int_pldif_8g_pld_tx_clk),
	.detectrxloopin(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdetectrxloopback),
	.dis_pc_byte(w_hssi_8g_rx_pcs_dis_pc_byte),
	.en_rev_parallel_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
	.hrdrst(gnd),
	.pcs_rst(\w_hssi_common_pcs_pma_interface_int_pmaif_8g_asn_bundling_in[3] ),
	.ph_fifo_rd_disable(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rddisable_tx),
	.pipe_en_rev_parallel_lpbk_in(w_hssi_tx_pld_pcs_interface_int_pldif_8g_rev_loopbk),
	.pipe_tx_deemph(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txdeemph),
	.rate_switch(w_hssi_8g_rx_pcs_gen2ngen1),
	.rd_enable_in_chnl_down(gnd),
	.rd_enable_in_chnl_up(gnd),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_8g_refclk_dig),
	.reset_pc_ptrs(w_hssi_8g_rx_pcs_reset_pc_ptrs),
	.reset_pc_ptrs_in_chnl_down(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_down_pipe),
	.reset_pc_ptrs_in_chnl_up(w_hssi_8g_rx_pcs_reset_pc_ptrs_in_chnl_up_pipe),
	.rxpolarity(w_hssi_rx_pld_pcs_interface_int_pldif_8g_rxpolarity),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_8g_scan_mode_n),
	.tx_pcs_reset(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txurstpcs_n),
	.txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
	.txswing(w_hssi_tx_pld_pcs_interface_int_pldif_8g_txswing),
	.wr_enable_in_chnl_down(gnd),
	.wr_enable_in_chnl_up(gnd),
	.wrenable_tx(w_hssi_tx_pld_pcs_interface_int_pldif_8g_wrenable_tx),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.bitslip_boundary_select({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[4] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[1] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_boundary_sel[0] }),
	.datain({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[40] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[39] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[36] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[34] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[32] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[29] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[28] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[20] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[19] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[16] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[14] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[12] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[9] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[8] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd[0] }),
	.eidleinfersel({\w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[2] ,\w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_8g_eidleinfersel[0] }),
	.fifo_select_in_chnl_down({gnd,gnd}),
	.fifo_select_in_chnl_up({gnd,gnd}),
	.pipe_tx_margin({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txmargin[0] }),
	.powerdn({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_powerdown[0] }),
	.rd_data_tx_phfifo({\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[63] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[62] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[61] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[60] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[59] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[58] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[57] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[56] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[55] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[54] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[53] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[52] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[51] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[50] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[49] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[48] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[47] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[46] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[45] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[44] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[43] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[42] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[41] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[40] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[39] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[38] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[37] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[36] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[35] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[34] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[33] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[32] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[31] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[30] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[29] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[28] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[27] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[26] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[25] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[24] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[23] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[22] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[21] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[20] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[19] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[18] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[17] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[16] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[15] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[14] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[13] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[12] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[11] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[10] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[9] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[8] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[7] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[6] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[5] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[4] ,
\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[3] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[2] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[1] ,\w_hssi_fifo_tx_pcs_data_out_8g_phase_comp[0] }),
	.rev_parallel_lpbk_data({\w_hssi_8g_rx_pcs_parallel_rev_loopback[19] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[18] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[17] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[16] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[15] ,
\w_hssi_8g_rx_pcs_parallel_rev_loopback[14] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[13] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[12] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[11] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[10] ,
\w_hssi_8g_rx_pcs_parallel_rev_loopback[9] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[8] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[7] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[6] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[5] ,
\w_hssi_8g_rx_pcs_parallel_rev_loopback[4] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[3] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[2] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[1] ,\w_hssi_8g_rx_pcs_parallel_rev_loopback[0] }),
	.tx_blk_start({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_blk_start[0] }),
	.tx_data_valid({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_data_valid[0] }),
	.tx_div_sync_in_chnl_down({gnd,gnd}),
	.tx_div_sync_in_chnl_up({gnd,gnd}),
	.tx_sync_hdr({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_tx_sync_hdr[0] }),
	.txd_fast_reg({\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[40] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[39] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[36] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[34] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[32] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[29] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[28] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[20] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[19] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[16] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[14] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[12] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[8] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_8g_txd_fast_reg[0] }),
	.blockselect(out_blockselect_hssi_8g_tx_pcs),
	.byte_serializer_pcs_clk_div_by_2_reg(),
	.byte_serializer_pcs_clk_div_by_2_wire(),
	.byte_serializer_pcs_clk_div_by_4_reg(),
	.byte_serializer_pld_clk_div_by_2_reg(),
	.byte_serializer_pld_clk_div_by_4_reg(),
	.clk_out(w_hssi_8g_tx_pcs_clk_out),
	.clk_out_gen3(w_hssi_8g_tx_pcs_clk_out_gen3),
	.dyn_clk_switch_n(w_hssi_8g_tx_pcs_dyn_clk_switch_n),
	.g3_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
	.g3_tx_pma_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
	.ph_fifo_overflow(w_hssi_8g_tx_pcs_ph_fifo_overflow),
	.ph_fifo_underflow(w_hssi_8g_tx_pcs_ph_fifo_underflow),
	.phfifo_txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
	.phfifo_txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
	.pipe_en_rev_parallel_lpbk_out(w_hssi_8g_tx_pcs_pipe_en_rev_parallel_lpbk_out),
	.pipe_tx_clk_out_gen3(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
	.pld_8g_empty_tx_fifo(),
	.pld_8g_empty_tx_reg(),
	.pld_8g_full_tx_fifo(),
	.pld_8g_full_tx_reg(),
	.pld_8g_g3_tx_pld_rst_n_reg(),
	.pld_8g_rddisable_tx_reg(),
	.pld_8g_tx_boundary_sel_reg(),
	.pld_pcs_tx_clk_out_8g_div_by_2_wire(),
	.pld_pcs_tx_clk_out_8g_wire(),
	.pld_tx_data_8g_fifo(),
	.pld_tx_data_lo_8g_reg(),
	.pmaif_asn_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
	.rd_enable_out_chnl_down(),
	.rd_enable_out_chnl_up(),
	.refclk_b(w_hssi_8g_tx_pcs_refclk_b),
	.refclk_b_reset(w_hssi_8g_tx_pcs_refclk_b_reset),
	.rxpolarity_int(w_hssi_8g_tx_pcs_rxpolarity_int),
	.soft_reset_wclk1_n(w_hssi_8g_tx_pcs_soft_reset_wclk1_n),
	.sta_tx_clk2_by2_1(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs~O_STA_TX_CLK2_BY2_1 ),
	.sta_tx_clk2_by2_1_out(),
	.sta_tx_clk2_by4_1(),
	.sta_tx_clk2_by4_1_out(),
	.sw_fifo_wr_clk(w_hssi_8g_tx_pcs_sw_fifo_wr_clk),
	.tx_clk_out_8g_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
	.tx_clk_out_pld_if(w_hssi_8g_tx_pcs_tx_clk_out_pld_if),
	.tx_clk_out_pmaif(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
	.tx_clk_to_observation_ff_in_pld_if(w_hssi_8g_tx_pcs_tx_clk_to_observation_ff_in_pld_if),
	.tx_detect_rxloopback_int(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
	.tx_pipe_clk(w_hssi_8g_tx_pcs_tx_pipe_clk),
	.tx_pipe_electidle(w_hssi_8g_tx_pcs_tx_pipe_electidle),
	.tx_pipe_soft_reset(w_hssi_8g_tx_pcs_tx_pipe_soft_reset),
	.txcompliance_out(w_hssi_8g_tx_pcs_txcompliance_out),
	.txelecidle_out(w_hssi_8g_tx_pcs_txelecidle_out),
	.wr_clk_tx_phfifo_dw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
	.wr_clk_tx_phfifo_sw_clk(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
	.wr_en_tx_phfifo(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
	.wr_enable_out_chnl_down(),
	.wr_enable_out_chnl_up(),
	.wr_rst_n_tx_phfifo(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
	.avmmreaddata(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_AVMMREADDATA_bus ),
	.dataout(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_DATAOUT_bus ),
	.fifo_select_out_chnl_down(),
	.fifo_select_out_chnl_up(),
	.non_gray_eidleinfersel(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_NON_GRAY_EIDLEINFERSEL_bus ),
	.phfifo_txmargin(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PHFIFO_TXMARGIN_bus ),
	.pipe_power_down_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_PIPE_POWER_DOWN_OUT_bus ),
	.rd_ptr_tx_phfifo(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_RD_PTR_TX_PHFIFO_bus ),
	.tx_blk_start_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_BLK_START_OUT_bus ),
	.tx_ctrlplane_testbus(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_CTRLPLANE_TESTBUS_bus ),
	.tx_data_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_OUT_bus ),
	.tx_data_valid_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATA_VALID_OUT_bus ),
	.tx_datak_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DATAK_OUT_bus ),
	.tx_div_sync(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_DIV_SYNC_bus ),
	.tx_div_sync_out_chnl_down(),
	.tx_div_sync_out_chnl_up(),
	.tx_sync_hdr_out(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_SYNC_HDR_OUT_bus ),
	.tx_testbus(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_TX_TESTBUS_bus ),
	.wr_data_tx_phfifo(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_DATA_TX_PHFIFO_bus ),
	.wr_ptr_tx_phfifo(\gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs_WR_PTR_TX_PHFIFO_bus ));
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .auto_speed_nego_gen2 = "dis_asn_g2";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .bit_reversal = "dis_bit_reversal";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .bonding_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .bonding_dft_val = "dft_0";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .bypass_pipeline_reg = "dis_bypass_pipeline";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .byte_serializer = "dis_bs";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .clock_gate_bs_enc = "dis_bs_enc_clk_gating";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .clock_gate_dw_fifowr = "en_dw_fifowr_clk_gating";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .clock_gate_fiford = "dis_fiford_clk_gating";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .clock_gate_sw_fifowr = "en_sw_fifowr_clk_gating";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .clock_observation_in_pld_core = "internal_refclk_b";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .ctrl_plane_bonding_compensation = "dis_compensation";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .ctrl_plane_bonding_consumption = "individual";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .ctrl_plane_bonding_distribution = "not_master_chnl_distr";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .data_selection_8b10b_encoder_input = "normal_data_path";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .dynamic_clk_switch = "dis_dyn_clk_switch";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .eightb_tenb_disp_ctrl = "dis_disp_ctrl";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .eightb_tenb_encoder = "en_8b10b_ibm";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .force_echar = "dis_force_echar";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .force_kchar = "dis_force_kchar";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .gen3_tx_clk_sel = "dis_tx_clk";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .gen3_tx_pipe_clk_sel = "dis_tx_pipe_clk";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .hip_mode = "dis_hip";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .pcs_bypass = "dis_pcs_bypass";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .phase_comp_rdptr = "disable_rdptr";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .phase_compensation_fifo = "register_fifo";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .phfifo_write_clk_sel = "tx_clk";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .pma_dw = "ten_bit";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .prot_mode = "cpri_rx_tx";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .refclk_b_clk_sel = "tx_pma_clock";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .revloop_back_rm = "dis_rev_loopback_rx_rm";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .symbol_swap = "dis_symbol_swap";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .tx_bitslip = "dis_tx_bitslip";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .tx_compliance_controlled_disparity = "dis_txcompliance";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .tx_fast_pld_reg = "dis_tx_fast_pld_reg";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .txclk_freerun = "en_freerun_tx";
defparam \gen_twentynm_hssi_8g_tx_pcs.inst_twentynm_hssi_8g_tx_pcs .txpcs_urst = "en_txpcs_urst";

twentynm_hssi_10g_tx_pcs \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.distdwn_in_dv(gnd),
	.distdwn_in_rden(gnd),
	.distdwn_in_wren(gnd),
	.distup_in_dv(gnd),
	.distup_in_rden(gnd),
	.distup_in_wren(gnd),
	.krfec_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_krfec_refclk_dig),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_10g_refclk_dig),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_10g_scan_mode_n),
	.tx_burst_en(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_burst_en),
	.tx_data_valid(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid),
	.tx_data_valid_reg(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_valid_reg),
	.tx_pld_clk(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_clk),
	.tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_pld_rst_n),
	.tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
	.tx_wordslip(w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_wordslip),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.r_tx_diag_word({gnd,vcc,vcc,gnd,gnd,vcc,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.r_tx_scrm_word({gnd,gnd,vcc,gnd,vcc,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.r_tx_skip_word({gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd}),
	.r_tx_sync_word({gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd,gnd,vcc,vcc,vcc,vcc,gnd,gnd,gnd,vcc,vcc,vcc,vcc,gnd,vcc,vcc,gnd}),
	.tx_bitslip({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[4] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[3] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_bitslip[0] }),
	.tx_control({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[16] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[14] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[12] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[10] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[8] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[6] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[4] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[2] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control[0] }),
	.tx_control_reg({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[8] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[5] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[4] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[1] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_control_reg[0] }),
	.tx_data({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[127] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[126] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[125] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[124] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[123] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[122] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[121] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[120] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[119] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[118] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[117] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[116] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[115] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[114] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[113] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[112] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[111] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[110] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[109] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[108] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[107] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[106] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[105] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[104] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[103] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[102] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[101] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[100] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[99] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[98] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[97] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[96] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[95] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[94] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[93] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[92] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[91] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[90] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[89] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[88] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[87] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[86] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[85] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[84] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[83] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[82] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[81] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[80] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[79] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[78] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[77] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[76] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[75] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[74] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[73] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[72] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[71] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[70] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[69] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[68] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[67] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[66] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[65] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[64] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[63] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[62] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[61] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[60] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[59] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[58] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[57] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[56] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[55] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[54] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[53] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[52] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[51] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[50] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[49] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[48] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[47] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[46] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[45] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[44] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[40] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[39] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[36] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[34] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[32] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[29] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[28] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[20] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[19] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[16] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[14] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[12] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[8] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data[0] }),
	.tx_data_in_krfec({\w_hssi_krfec_tx_pcs_tx_data_out[63] ,\w_hssi_krfec_tx_pcs_tx_data_out[62] ,\w_hssi_krfec_tx_pcs_tx_data_out[61] ,\w_hssi_krfec_tx_pcs_tx_data_out[60] ,\w_hssi_krfec_tx_pcs_tx_data_out[59] ,\w_hssi_krfec_tx_pcs_tx_data_out[58] ,
\w_hssi_krfec_tx_pcs_tx_data_out[57] ,\w_hssi_krfec_tx_pcs_tx_data_out[56] ,\w_hssi_krfec_tx_pcs_tx_data_out[55] ,\w_hssi_krfec_tx_pcs_tx_data_out[54] ,\w_hssi_krfec_tx_pcs_tx_data_out[53] ,\w_hssi_krfec_tx_pcs_tx_data_out[52] ,
\w_hssi_krfec_tx_pcs_tx_data_out[51] ,\w_hssi_krfec_tx_pcs_tx_data_out[50] ,\w_hssi_krfec_tx_pcs_tx_data_out[49] ,\w_hssi_krfec_tx_pcs_tx_data_out[48] ,\w_hssi_krfec_tx_pcs_tx_data_out[47] ,\w_hssi_krfec_tx_pcs_tx_data_out[46] ,
\w_hssi_krfec_tx_pcs_tx_data_out[45] ,\w_hssi_krfec_tx_pcs_tx_data_out[44] ,\w_hssi_krfec_tx_pcs_tx_data_out[43] ,\w_hssi_krfec_tx_pcs_tx_data_out[42] ,\w_hssi_krfec_tx_pcs_tx_data_out[41] ,\w_hssi_krfec_tx_pcs_tx_data_out[40] ,
\w_hssi_krfec_tx_pcs_tx_data_out[39] ,\w_hssi_krfec_tx_pcs_tx_data_out[38] ,\w_hssi_krfec_tx_pcs_tx_data_out[37] ,\w_hssi_krfec_tx_pcs_tx_data_out[36] ,\w_hssi_krfec_tx_pcs_tx_data_out[35] ,\w_hssi_krfec_tx_pcs_tx_data_out[34] ,
\w_hssi_krfec_tx_pcs_tx_data_out[33] ,\w_hssi_krfec_tx_pcs_tx_data_out[32] ,\w_hssi_krfec_tx_pcs_tx_data_out[31] ,\w_hssi_krfec_tx_pcs_tx_data_out[30] ,\w_hssi_krfec_tx_pcs_tx_data_out[29] ,\w_hssi_krfec_tx_pcs_tx_data_out[28] ,
\w_hssi_krfec_tx_pcs_tx_data_out[27] ,\w_hssi_krfec_tx_pcs_tx_data_out[26] ,\w_hssi_krfec_tx_pcs_tx_data_out[25] ,\w_hssi_krfec_tx_pcs_tx_data_out[24] ,\w_hssi_krfec_tx_pcs_tx_data_out[23] ,\w_hssi_krfec_tx_pcs_tx_data_out[22] ,
\w_hssi_krfec_tx_pcs_tx_data_out[21] ,\w_hssi_krfec_tx_pcs_tx_data_out[20] ,\w_hssi_krfec_tx_pcs_tx_data_out[19] ,\w_hssi_krfec_tx_pcs_tx_data_out[18] ,\w_hssi_krfec_tx_pcs_tx_data_out[17] ,\w_hssi_krfec_tx_pcs_tx_data_out[16] ,
\w_hssi_krfec_tx_pcs_tx_data_out[15] ,\w_hssi_krfec_tx_pcs_tx_data_out[14] ,\w_hssi_krfec_tx_pcs_tx_data_out[13] ,\w_hssi_krfec_tx_pcs_tx_data_out[12] ,\w_hssi_krfec_tx_pcs_tx_data_out[11] ,\w_hssi_krfec_tx_pcs_tx_data_out[10] ,
\w_hssi_krfec_tx_pcs_tx_data_out[9] ,\w_hssi_krfec_tx_pcs_tx_data_out[8] ,\w_hssi_krfec_tx_pcs_tx_data_out[7] ,\w_hssi_krfec_tx_pcs_tx_data_out[6] ,\w_hssi_krfec_tx_pcs_tx_data_out[5] ,\w_hssi_krfec_tx_pcs_tx_data_out[4] ,\w_hssi_krfec_tx_pcs_tx_data_out[3] ,
\w_hssi_krfec_tx_pcs_tx_data_out[2] ,\w_hssi_krfec_tx_pcs_tx_data_out[1] ,\w_hssi_krfec_tx_pcs_tx_data_out[0] }),
	.tx_data_reg({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[63] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[62] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[61] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[60] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[59] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[58] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[57] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[56] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[55] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[54] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[53] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[52] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[51] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[50] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[49] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[48] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[47] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[46] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[45] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[44] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[40] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[39] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[36] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[34] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[32] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[29] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[28] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[20] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[19] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[16] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[14] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[12] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[8] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_data_reg[0] }),
	.tx_diag_status({\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_10g_tx_diag_status[0] }),
	.tx_fifo_rd_data({\w_hssi_fifo_tx_pcs_data_out_10g[72] ,\w_hssi_fifo_tx_pcs_data_out_10g[71] ,\w_hssi_fifo_tx_pcs_data_out_10g[70] ,\w_hssi_fifo_tx_pcs_data_out_10g[69] ,\w_hssi_fifo_tx_pcs_data_out_10g[68] ,\w_hssi_fifo_tx_pcs_data_out_10g[67] ,
\w_hssi_fifo_tx_pcs_data_out_10g[66] ,\w_hssi_fifo_tx_pcs_data_out_10g[65] ,\w_hssi_fifo_tx_pcs_data_out_10g[64] ,\w_hssi_fifo_tx_pcs_data_out_10g[63] ,\w_hssi_fifo_tx_pcs_data_out_10g[62] ,\w_hssi_fifo_tx_pcs_data_out_10g[61] ,
\w_hssi_fifo_tx_pcs_data_out_10g[60] ,\w_hssi_fifo_tx_pcs_data_out_10g[59] ,\w_hssi_fifo_tx_pcs_data_out_10g[58] ,\w_hssi_fifo_tx_pcs_data_out_10g[57] ,\w_hssi_fifo_tx_pcs_data_out_10g[56] ,\w_hssi_fifo_tx_pcs_data_out_10g[55] ,
\w_hssi_fifo_tx_pcs_data_out_10g[54] ,\w_hssi_fifo_tx_pcs_data_out_10g[53] ,\w_hssi_fifo_tx_pcs_data_out_10g[52] ,\w_hssi_fifo_tx_pcs_data_out_10g[51] ,\w_hssi_fifo_tx_pcs_data_out_10g[50] ,\w_hssi_fifo_tx_pcs_data_out_10g[49] ,
\w_hssi_fifo_tx_pcs_data_out_10g[48] ,\w_hssi_fifo_tx_pcs_data_out_10g[47] ,\w_hssi_fifo_tx_pcs_data_out_10g[46] ,\w_hssi_fifo_tx_pcs_data_out_10g[45] ,\w_hssi_fifo_tx_pcs_data_out_10g[44] ,\w_hssi_fifo_tx_pcs_data_out_10g[43] ,
\w_hssi_fifo_tx_pcs_data_out_10g[42] ,\w_hssi_fifo_tx_pcs_data_out_10g[41] ,\w_hssi_fifo_tx_pcs_data_out_10g[40] ,\w_hssi_fifo_tx_pcs_data_out_10g[39] ,\w_hssi_fifo_tx_pcs_data_out_10g[38] ,\w_hssi_fifo_tx_pcs_data_out_10g[37] ,
\w_hssi_fifo_tx_pcs_data_out_10g[36] ,\w_hssi_fifo_tx_pcs_data_out_10g[35] ,\w_hssi_fifo_tx_pcs_data_out_10g[34] ,\w_hssi_fifo_tx_pcs_data_out_10g[33] ,\w_hssi_fifo_tx_pcs_data_out_10g[32] ,\w_hssi_fifo_tx_pcs_data_out_10g[31] ,
\w_hssi_fifo_tx_pcs_data_out_10g[30] ,\w_hssi_fifo_tx_pcs_data_out_10g[29] ,\w_hssi_fifo_tx_pcs_data_out_10g[28] ,\w_hssi_fifo_tx_pcs_data_out_10g[27] ,\w_hssi_fifo_tx_pcs_data_out_10g[26] ,\w_hssi_fifo_tx_pcs_data_out_10g[25] ,
\w_hssi_fifo_tx_pcs_data_out_10g[24] ,\w_hssi_fifo_tx_pcs_data_out_10g[23] ,\w_hssi_fifo_tx_pcs_data_out_10g[22] ,\w_hssi_fifo_tx_pcs_data_out_10g[21] ,\w_hssi_fifo_tx_pcs_data_out_10g[20] ,\w_hssi_fifo_tx_pcs_data_out_10g[19] ,
\w_hssi_fifo_tx_pcs_data_out_10g[18] ,\w_hssi_fifo_tx_pcs_data_out_10g[17] ,\w_hssi_fifo_tx_pcs_data_out_10g[16] ,\w_hssi_fifo_tx_pcs_data_out_10g[15] ,\w_hssi_fifo_tx_pcs_data_out_10g[14] ,\w_hssi_fifo_tx_pcs_data_out_10g[13] ,
\w_hssi_fifo_tx_pcs_data_out_10g[12] ,\w_hssi_fifo_tx_pcs_data_out_10g[11] ,\w_hssi_fifo_tx_pcs_data_out_10g[10] ,\w_hssi_fifo_tx_pcs_data_out_10g[9] ,\w_hssi_fifo_tx_pcs_data_out_10g[8] ,\w_hssi_fifo_tx_pcs_data_out_10g[7] ,\w_hssi_fifo_tx_pcs_data_out_10g[6] ,
\w_hssi_fifo_tx_pcs_data_out_10g[5] ,\w_hssi_fifo_tx_pcs_data_out_10g[4] ,\w_hssi_fifo_tx_pcs_data_out_10g[3] ,\w_hssi_fifo_tx_pcs_data_out_10g[2] ,\w_hssi_fifo_tx_pcs_data_out_10g[1] ,\w_hssi_fifo_tx_pcs_data_out_10g[0] }),
	.blockselect(out_blockselect_hssi_10g_tx_pcs),
	.distdwn_out_dv(),
	.distdwn_out_rden(),
	.distdwn_out_wren(),
	.distup_out_dv(),
	.distup_out_rden(),
	.distup_out_wren(),
	.pld_10g_krfec_tx_frame_10g_reg(),
	.pld_10g_krfec_tx_pld_rst_n_fifo(),
	.pld_10g_krfec_tx_pld_rst_n_reg(),
	.pld_10g_tx_bitslip_reg(),
	.pld_10g_tx_burst_en_exe_reg(),
	.pld_10g_tx_data_valid_10g_reg(),
	.pld_10g_tx_data_valid_fifo(),
	.pld_10g_tx_data_valid_reg(),
	.pld_10g_tx_diag_status_reg(),
	.pld_10g_tx_empty_reg(),
	.pld_10g_tx_fifo_num_reg(),
	.pld_10g_tx_full_fifo(),
	.pld_10g_tx_full_reg(),
	.pld_10g_tx_pempty_reg(),
	.pld_10g_tx_pfull_fifo(),
	.pld_10g_tx_wordslip_exe_reg(),
	.pld_10g_tx_wordslip_reg(),
	.pld_pcs_tx_clk_out_10g_wire(),
	.pld_tx_burst_en_reg(),
	.pld_tx_control_lo_10g_reg(),
	.pld_tx_data_10g_fifo(),
	.pld_tx_data_lo_10g_reg(),
	.tx_burst_en_exe(w_hssi_10g_tx_pcs_tx_burst_en_exe),
	.tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out),
	.tx_clk_out_pld_if(w_hssi_10g_tx_pcs_tx_clk_out_pld_if),
	.tx_clk_out_pma_if(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
	.tx_data_valid_out_krfec(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
	.tx_dft_clk_out(w_hssi_10g_tx_pcs_tx_dft_clk_out),
	.tx_empty(w_hssi_10g_tx_pcs_tx_empty),
	.tx_fec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
	.tx_fifo_wr_clk(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
	.tx_fifo_wr_en(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
	.tx_fifo_wr_rst_n(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
	.tx_frame(w_hssi_10g_tx_pcs_tx_frame),
	.tx_full(w_hssi_10g_tx_pcs_tx_full),
	.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
	.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
	.tx_pempty(w_hssi_10g_tx_pcs_tx_pempty),
	.tx_pfull(w_hssi_10g_tx_pcs_tx_pfull),
	.tx_wordslip_exe(w_hssi_10g_tx_pcs_tx_wordslip_exe),
	.avmmreaddata(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_AVMMREADDATA_bus ),
	.tx_control_out_krfec(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_CONTROL_OUT_KRFEC_bus ),
	.tx_data_out_krfec(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_DATA_OUT_KRFEC_bus ),
	.tx_fifo_num(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_NUM_bus ),
	.tx_fifo_rd_ptr(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_RD_PTR_bus ),
	.tx_fifo_wr_data(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_bus ),
	.tx_fifo_wr_data_dw(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_DATA_DW_bus ),
	.tx_fifo_wr_ptr(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_FIFO_WR_PTR_bus ),
	.tx_pma_data(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_DATA_bus ),
	.tx_pma_gating_val(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_PMA_GATING_VAL_bus ),
	.tx_test_data(\gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs_TX_TEST_DATA_bus ));
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .advanced_user_mode = "disable";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .bitslip_en = "bitslip_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .bonding_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .bonding_dft_val = "dft_0";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .comp_cnt = 8'b00000000;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .compin_sel = "compin_master";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .crcgen_bypass = "crcgen_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .crcgen_clken = "crcgen_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .crcgen_err = "crcgen_err_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .crcgen_inv = "crcgen_inv_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .ctrl_bit_reverse = "ctrl_bit_reverse_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .ctrl_plane_bonding = "individual";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .data_bit_reverse = "data_bit_reverse_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dft_clk_out_sel = "tx_master_clk";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dispgen_bypass = "dispgen_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dispgen_clken = "dispgen_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dispgen_err = "dispgen_err_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dispgen_pipeln = "dispgen_pipeln_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .distdwn_bypass_pipeln = "distdwn_bypass_pipeln_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .distdwn_master = "distdwn_master_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .distup_bypass_pipeln = "distup_bypass_pipeln_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .distup_master = "distup_master_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .dv_bond = "dv_bond_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .empty_flag_type = "empty_rd_side";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .enc64b66b_txsm_clken = "enc64b66b_txsm_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .enc_64b66b_txsm_bypass = "enc_64b66b_txsm_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fastpath = "fastpath_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fec_clken = "fec_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fec_enable = "fec_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fifo_double_write = "fifo_double_write_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fifo_reg_fast = "fifo_reg_fast_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fifo_stop_rd = "rd_empty";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .fifo_stop_wr = "n_wr_full";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_burst = "frmgen_burst_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_bypass = "frmgen_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_clken = "frmgen_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_mfrm_length = 16'b0000100000000000;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_pipeln = "frmgen_pipeln_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_pyld_ins = "frmgen_pyld_ins_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .frmgen_wordslip = "frmgen_wordslip_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .full_flag_type = "full_wr_side";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .gb_pipeln_bypass = "disable";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .gb_tx_idwidth = "width_64";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .gb_tx_odwidth = "width_64";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .gbred_clken = "gbred_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .indv = "indv_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .low_latency_en = "disable";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .master_clk_sel = "master_tx_pma_clk";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pempty_flag_type = "pempty_rd_side";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pfull_flag_type = "pfull_wr_side";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .phcomp_rd_del = "phcomp_rd_del2";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pld_if_type = "fifo";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .prot_mode = "disable_mode";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pseudo_random = "all_0";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pseudo_seed_a = 58'b1111111111111111111111111111111111111111111111111111111111;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .pseudo_seed_b = 58'b1111111111111111111111111111111111111111111111111111111111;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .random_disp = "disable";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .rdfifo_clken = "rdfifo_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .scrm_bypass = "scrm_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .scrm_clken = "scrm_clk_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .scrm_mode = "async";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .scrm_pipeln = "enable";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .sh_err = "sh_err_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .sop_mark = "sop_mark_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .stretch_num_stages = "zero_stage";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .test_mode = "test_off";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_scrm_err = "scrm_err_dis";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_scrm_width = "bit64";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_sh_location = "msb";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_sm_bypass = "tx_sm_bypass_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_sm_pipeln = "tx_sm_pipeln_en";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .tx_testbus_sel = "tx_fifo_testbus1";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .txfifo_empty = "empty_default";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .txfifo_full = "full_default";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .txfifo_mode = "phase_comp";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .txfifo_pempty = 4'b0010;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .txfifo_pfull = 4'b1011;
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .wr_clk_sel = "wr_tx_pld_clk";
defparam \gen_twentynm_hssi_10g_tx_pcs.inst_twentynm_hssi_10g_tx_pcs .wrfifo_clken = "wrfifo_clk_dis";

twentynm_hssi_gen3_rx_pcs \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
	.inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
	.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
	.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
	.rcvd_clk(w_hssi_8g_rx_pcs_rx_rcvd_clk_gen3),
	.rx_pma_clk(w_hssi_8g_rx_pcs_rx_pma_clk_gen3),
	.rx_pma_rstn(w_hssi_8g_rx_pcs_g3_rx_pma_rstn),
	.rx_rcvd_rstn(w_hssi_8g_rx_pcs_g3_rx_rcvd_rstn),
	.rxpolarity(w_hssi_pipe_gen3_rxpolarity_int),
	.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
	.sync_sm_en(w_hssi_rx_pld_pcs_interface_int_pldif_g3_syncsm_en),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.data_in({\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[31] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[30] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[29] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[28] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[27] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[26] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[25] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[24] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[23] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[22] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[21] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[20] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[19] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[18] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[17] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[16] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[15] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[14] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[13] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[12] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[11] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[10] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[9] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[8] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[7] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[6] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[5] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[4] ,
\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[3] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[2] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[1] ,\w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_data_in[0] }),
	.mem_rx_fifo_rd_data({\w_hssi_fifo_rx_pcs_data_out_gen3[39] ,\w_hssi_fifo_rx_pcs_data_out_gen3[38] ,\w_hssi_fifo_rx_pcs_data_out_gen3[37] ,\w_hssi_fifo_rx_pcs_data_out_gen3[36] ,\w_hssi_fifo_rx_pcs_data_out_gen3[35] ,\w_hssi_fifo_rx_pcs_data_out_gen3[34] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[33] ,\w_hssi_fifo_rx_pcs_data_out_gen3[32] ,\w_hssi_fifo_rx_pcs_data_out_gen3[31] ,\w_hssi_fifo_rx_pcs_data_out_gen3[30] ,\w_hssi_fifo_rx_pcs_data_out_gen3[29] ,\w_hssi_fifo_rx_pcs_data_out_gen3[28] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[27] ,\w_hssi_fifo_rx_pcs_data_out_gen3[26] ,\w_hssi_fifo_rx_pcs_data_out_gen3[25] ,\w_hssi_fifo_rx_pcs_data_out_gen3[24] ,\w_hssi_fifo_rx_pcs_data_out_gen3[23] ,\w_hssi_fifo_rx_pcs_data_out_gen3[22] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[21] ,\w_hssi_fifo_rx_pcs_data_out_gen3[20] ,\w_hssi_fifo_rx_pcs_data_out_gen3[19] ,\w_hssi_fifo_rx_pcs_data_out_gen3[18] ,\w_hssi_fifo_rx_pcs_data_out_gen3[17] ,\w_hssi_fifo_rx_pcs_data_out_gen3[16] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[15] ,\w_hssi_fifo_rx_pcs_data_out_gen3[14] ,\w_hssi_fifo_rx_pcs_data_out_gen3[13] ,\w_hssi_fifo_rx_pcs_data_out_gen3[12] ,\w_hssi_fifo_rx_pcs_data_out_gen3[11] ,\w_hssi_fifo_rx_pcs_data_out_gen3[10] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[9] ,\w_hssi_fifo_rx_pcs_data_out_gen3[8] ,\w_hssi_fifo_rx_pcs_data_out_gen3[7] ,\w_hssi_fifo_rx_pcs_data_out_gen3[6] ,\w_hssi_fifo_rx_pcs_data_out_gen3[5] ,\w_hssi_fifo_rx_pcs_data_out_gen3[4] ,
\w_hssi_fifo_rx_pcs_data_out_gen3[3] ,\w_hssi_fifo_rx_pcs_data_out_gen3[2] ,\w_hssi_fifo_rx_pcs_data_out_gen3[1] ,\w_hssi_fifo_rx_pcs_data_out_gen3[0] }),
	.par_lpbk_b4gb_in({\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[35] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[34] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[33] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[32] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[31] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[30] ,
\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[29] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[28] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[27] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[26] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[25] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[24] ,
\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[23] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[22] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[21] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[20] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[19] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[18] ,
\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[17] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[16] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[15] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[14] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[13] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[12] ,
\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[11] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[10] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[9] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[8] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[7] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[6] ,
\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[5] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[4] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[3] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[2] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[1] ,\w_hssi_gen3_tx_pcs_par_lpbk_b4gb_out[0] }),
	.par_lpbk_in({\w_hssi_gen3_tx_pcs_par_lpbk_out[31] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[30] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[29] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[28] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[27] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[26] ,
\w_hssi_gen3_tx_pcs_par_lpbk_out[25] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[24] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[23] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[22] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[21] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[20] ,
\w_hssi_gen3_tx_pcs_par_lpbk_out[19] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[18] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[17] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[16] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[15] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[14] ,
\w_hssi_gen3_tx_pcs_par_lpbk_out[13] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[12] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[11] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[10] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[9] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[8] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[7] ,
\w_hssi_gen3_tx_pcs_par_lpbk_out[6] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[5] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[4] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[3] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[2] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[1] ,\w_hssi_gen3_tx_pcs_par_lpbk_out[0] }),
	.txdatak_in({\w_hssi_pipe_gen3_txdatak_int[3] ,\w_hssi_pipe_gen3_txdatak_int[2] ,\w_hssi_pipe_gen3_txdatak_int[1] ,\w_hssi_pipe_gen3_txdatak_int[0] }),
	.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
	.blk_lockd_int(),
	.blk_start(w_hssi_gen3_rx_pcs_blk_start),
	.blockselect(out_blockselect_hssi_gen3_rx_pcs),
	.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
	.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
	.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
	.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
	.data_valid(w_hssi_gen3_rx_pcs_data_valid),
	.ei_det_int(w_hssi_gen3_rx_pcs_ei_det_int),
	.ei_partial_det_int(w_hssi_gen3_rx_pcs_ei_partial_det_int),
	.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
	.i_det_int(w_hssi_gen3_rx_pcs_i_det_int),
	.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
	.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
	.mem_rx_fifo_wr_clk(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
	.mem_rx_fifo_wr_en(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
	.mem_rx_fifo_wr_rst_n(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
	.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
	.skp_det_int(),
	.avmmreaddata(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_AVMMREADDATA_bus ),
	.data_out(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_DATA_OUT_bus ),
	.lpbk_data(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_LPBK_DATA_bus ),
	.mem_rx_fifo_rd_ptr(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_RD_PTR_bus ),
	.mem_rx_fifo_wr_data(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_DATA_bus ),
	.mem_rx_fifo_wr_ptr(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_MEM_RX_FIFO_WR_PTR_bus ),
	.rx_test_out(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_RX_TEST_OUT_bus ),
	.sync_hdr(\gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs_SYNC_HDR_bus ));
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .block_sync = "bypass_block_sync";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .block_sync_sm = "disable_blk_sync_sm";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .cdr_ctrl_force_unalgn = "disable";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .lpbk_force = "lpbk_frce_dis";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .mode = "disable_pcs";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rate_match_fifo = "bypass_rm_fifo";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rate_match_fifo_latency = "low_latency";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .reverse_lpbk = "rev_lpbk_dis";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rx_b4gb_par_lpbk = "b4gb_par_lpbk_dis";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rx_force_balign = "dis_force_balign";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rx_ins_del_one_skip = "ins_del_one_skip_dis";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rx_num_fixed_pat = 4'b0000;
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .rx_test_out_sel = "rx_test_out0";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_gen3_rx_pcs.inst_twentynm_hssi_gen3_rx_pcs .sup_mode = "user_mode";

twentynm_hssi_pipe_gen3 \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.blk_algnd_int(w_hssi_gen3_rx_pcs_blk_algnd_int),
	.clkcomp_delete_int(w_hssi_gen3_rx_pcs_clkcomp_delete_int),
	.clkcomp_insert_int(w_hssi_gen3_rx_pcs_clkcomp_insert_int),
	.clkcomp_overfl_int(w_hssi_gen3_rx_pcs_clkcomp_overfl_int),
	.clkcomp_undfl_int(w_hssi_gen3_rx_pcs_clkcomp_undfl_int),
	.err_decode_int(w_hssi_gen3_rx_pcs_err_decode_int),
	.pipe_tx_clk(w_hssi_8g_tx_pcs_pipe_tx_clk_out_gen3),
	.pipe_tx_rstn(w_hssi_8g_tx_pcs_g3_pipe_tx_pma_rstn),
	.pma_rx_detect_valid(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_detect_valid),
	.pma_rx_found(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_rx_found),
	.pma_signal_det(w_hssi_rx_pcs_pma_interface_int_pmaif_g3_pma_signal_det),
	.rcv_lfsr_chk_int(w_hssi_gen3_rx_pcs_rcv_lfsr_chk_int),
	.rx_blk_start_int(w_hssi_gen3_rx_pcs_blk_start),
	.rxdataskip_int(w_hssi_gen3_rx_pcs_data_valid),
	.rxelecidle_8gpcs_in(w_hssi_pipe_gen1_2_rxelectricalidle_out),
	.rxpolarity(w_hssi_8g_tx_pcs_rxpolarity_int),
	.tx_blk_start(\w_hssi_8g_tx_pcs_tx_blk_start_out[0] ),
	.txcompliance(w_hssi_8g_tx_pcs_txcompliance_out),
	.txdataskip(\w_hssi_8g_tx_pcs_tx_data_valid_out[0] ),
	.txdeemph(w_hssi_8g_tx_pcs_phfifo_txdeemph),
	.txdetectrxloopback(w_hssi_8g_tx_pcs_tx_detect_rxloopback_int),
	.txelecidle(w_hssi_8g_tx_pcs_txelecidle_out),
	.txswing(w_hssi_8g_tx_pcs_phfifo_txswing),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.current_coeff({\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[17] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[16] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[15] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[14] ,
\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[13] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[12] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[11] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[10] ,
\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[9] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[8] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[7] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[6] ,
\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[5] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[4] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[3] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[2] ,
\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_coeff[0] }),
	.current_rxpreset({\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[2] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_g3_current_rxpreset[0] }),
	.pcs_asn_bundling_in({\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[8] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[7] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[6] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[5] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[4] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[3] ,
\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[2] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[1] ,\w_hssi_common_pcs_pma_interface_int_pmaif_g3_pcs_asn_bundling_in[0] }),
	.powerdown({\w_hssi_8g_tx_pcs_pipe_power_down_out[1] ,\w_hssi_8g_tx_pcs_pipe_power_down_out[0] }),
	.rx_sync_hdr_int({\w_hssi_gen3_rx_pcs_sync_hdr[1] ,\w_hssi_gen3_rx_pcs_sync_hdr[0] }),
	.rx_test_out({\w_hssi_gen3_rx_pcs_rx_test_out[19] ,\w_hssi_gen3_rx_pcs_rx_test_out[18] ,\w_hssi_gen3_rx_pcs_rx_test_out[17] ,\w_hssi_gen3_rx_pcs_rx_test_out[16] ,\w_hssi_gen3_rx_pcs_rx_test_out[15] ,\w_hssi_gen3_rx_pcs_rx_test_out[14] ,\w_hssi_gen3_rx_pcs_rx_test_out[13] ,
\w_hssi_gen3_rx_pcs_rx_test_out[12] ,\w_hssi_gen3_rx_pcs_rx_test_out[11] ,\w_hssi_gen3_rx_pcs_rx_test_out[10] ,\w_hssi_gen3_rx_pcs_rx_test_out[9] ,\w_hssi_gen3_rx_pcs_rx_test_out[8] ,\w_hssi_gen3_rx_pcs_rx_test_out[7] ,\w_hssi_gen3_rx_pcs_rx_test_out[6] ,
\w_hssi_gen3_rx_pcs_rx_test_out[5] ,\w_hssi_gen3_rx_pcs_rx_test_out[4] ,\w_hssi_gen3_rx_pcs_rx_test_out[3] ,\w_hssi_gen3_rx_pcs_rx_test_out[2] ,\w_hssi_gen3_rx_pcs_rx_test_out[1] ,\w_hssi_gen3_rx_pcs_rx_test_out[0] }),
	.rxd_8gpcs_in({\w_hssi_8g_rx_pcs_pipe_data[63] ,\w_hssi_8g_rx_pcs_pipe_data[62] ,\w_hssi_8g_rx_pcs_pipe_data[61] ,\w_hssi_8g_rx_pcs_pipe_data[60] ,\w_hssi_8g_rx_pcs_pipe_data[59] ,\w_hssi_8g_rx_pcs_pipe_data[58] ,\w_hssi_8g_rx_pcs_pipe_data[57] ,\w_hssi_8g_rx_pcs_pipe_data[56] ,
\w_hssi_8g_rx_pcs_pipe_data[55] ,\w_hssi_8g_rx_pcs_pipe_data[54] ,\w_hssi_8g_rx_pcs_pipe_data[53] ,\w_hssi_8g_rx_pcs_pipe_data[52] ,\w_hssi_8g_rx_pcs_pipe_data[51] ,\w_hssi_8g_rx_pcs_pipe_data[50] ,\w_hssi_8g_rx_pcs_pipe_data[49] ,\w_hssi_8g_rx_pcs_pipe_data[48] ,
\w_hssi_8g_rx_pcs_pipe_data[47] ,\w_hssi_8g_rx_pcs_pipe_data[46] ,\w_hssi_8g_rx_pcs_pipe_data[45] ,\w_hssi_8g_rx_pcs_pipe_data[44] ,\w_hssi_8g_rx_pcs_pipe_data[43] ,\w_hssi_8g_rx_pcs_pipe_data[42] ,\w_hssi_8g_rx_pcs_pipe_data[41] ,\w_hssi_8g_rx_pcs_pipe_data[40] ,
\w_hssi_8g_rx_pcs_pipe_data[39] ,\w_hssi_8g_rx_pcs_pipe_data[38] ,\w_hssi_8g_rx_pcs_pipe_data[37] ,\w_hssi_8g_rx_pcs_pipe_data[36] ,\w_hssi_8g_rx_pcs_pipe_data[35] ,\w_hssi_8g_rx_pcs_pipe_data[34] ,\w_hssi_8g_rx_pcs_pipe_data[33] ,\w_hssi_8g_rx_pcs_pipe_data[32] ,
\w_hssi_8g_rx_pcs_pipe_data[31] ,\w_hssi_8g_rx_pcs_pipe_data[30] ,\w_hssi_8g_rx_pcs_pipe_data[29] ,\w_hssi_8g_rx_pcs_pipe_data[28] ,\w_hssi_8g_rx_pcs_pipe_data[27] ,\w_hssi_8g_rx_pcs_pipe_data[26] ,\w_hssi_8g_rx_pcs_pipe_data[25] ,\w_hssi_8g_rx_pcs_pipe_data[24] ,
\w_hssi_8g_rx_pcs_pipe_data[23] ,\w_hssi_8g_rx_pcs_pipe_data[22] ,\w_hssi_8g_rx_pcs_pipe_data[21] ,\w_hssi_8g_rx_pcs_pipe_data[20] ,\w_hssi_8g_rx_pcs_pipe_data[19] ,\w_hssi_8g_rx_pcs_pipe_data[18] ,\w_hssi_8g_rx_pcs_pipe_data[17] ,\w_hssi_8g_rx_pcs_pipe_data[16] ,
\w_hssi_8g_rx_pcs_pipe_data[15] ,\w_hssi_8g_rx_pcs_pipe_data[14] ,\w_hssi_8g_rx_pcs_pipe_data[13] ,\w_hssi_8g_rx_pcs_pipe_data[12] ,\w_hssi_8g_rx_pcs_pipe_data[11] ,\w_hssi_8g_rx_pcs_pipe_data[10] ,\w_hssi_8g_rx_pcs_pipe_data[9] ,\w_hssi_8g_rx_pcs_pipe_data[8] ,
\w_hssi_8g_rx_pcs_pipe_data[7] ,\w_hssi_8g_rx_pcs_pipe_data[6] ,\w_hssi_8g_rx_pcs_pipe_data[5] ,\w_hssi_8g_rx_pcs_pipe_data[4] ,\w_hssi_8g_rx_pcs_pipe_data[3] ,\w_hssi_8g_rx_pcs_pipe_data[2] ,\w_hssi_8g_rx_pcs_pipe_data[1] ,\w_hssi_8g_rx_pcs_pipe_data[0] }),
	.rxdata_int({\w_hssi_gen3_rx_pcs_data_out[31] ,\w_hssi_gen3_rx_pcs_data_out[30] ,\w_hssi_gen3_rx_pcs_data_out[29] ,\w_hssi_gen3_rx_pcs_data_out[28] ,\w_hssi_gen3_rx_pcs_data_out[27] ,\w_hssi_gen3_rx_pcs_data_out[26] ,\w_hssi_gen3_rx_pcs_data_out[25] ,
\w_hssi_gen3_rx_pcs_data_out[24] ,\w_hssi_gen3_rx_pcs_data_out[23] ,\w_hssi_gen3_rx_pcs_data_out[22] ,\w_hssi_gen3_rx_pcs_data_out[21] ,\w_hssi_gen3_rx_pcs_data_out[20] ,\w_hssi_gen3_rx_pcs_data_out[19] ,\w_hssi_gen3_rx_pcs_data_out[18] ,
\w_hssi_gen3_rx_pcs_data_out[17] ,\w_hssi_gen3_rx_pcs_data_out[16] ,\w_hssi_gen3_rx_pcs_data_out[15] ,\w_hssi_gen3_rx_pcs_data_out[14] ,\w_hssi_gen3_rx_pcs_data_out[13] ,\w_hssi_gen3_rx_pcs_data_out[12] ,\w_hssi_gen3_rx_pcs_data_out[11] ,
\w_hssi_gen3_rx_pcs_data_out[10] ,\w_hssi_gen3_rx_pcs_data_out[9] ,\w_hssi_gen3_rx_pcs_data_out[8] ,\w_hssi_gen3_rx_pcs_data_out[7] ,\w_hssi_gen3_rx_pcs_data_out[6] ,\w_hssi_gen3_rx_pcs_data_out[5] ,\w_hssi_gen3_rx_pcs_data_out[4] ,
\w_hssi_gen3_rx_pcs_data_out[3] ,\w_hssi_gen3_rx_pcs_data_out[2] ,\w_hssi_gen3_rx_pcs_data_out[1] ,\w_hssi_gen3_rx_pcs_data_out[0] }),
	.rxdatak_int({gnd,gnd,gnd,gnd}),
	.tx_sync_hdr({\w_hssi_8g_tx_pcs_tx_sync_hdr_out[1] ,\w_hssi_8g_tx_pcs_tx_sync_hdr_out[0] }),
	.tx_test_out({\w_hssi_gen3_tx_pcs_tx_test_out[19] ,\w_hssi_gen3_tx_pcs_tx_test_out[18] ,\w_hssi_gen3_tx_pcs_tx_test_out[17] ,\w_hssi_gen3_tx_pcs_tx_test_out[16] ,\w_hssi_gen3_tx_pcs_tx_test_out[15] ,\w_hssi_gen3_tx_pcs_tx_test_out[14] ,\w_hssi_gen3_tx_pcs_tx_test_out[13] ,
\w_hssi_gen3_tx_pcs_tx_test_out[12] ,\w_hssi_gen3_tx_pcs_tx_test_out[11] ,\w_hssi_gen3_tx_pcs_tx_test_out[10] ,\w_hssi_gen3_tx_pcs_tx_test_out[9] ,\w_hssi_gen3_tx_pcs_tx_test_out[8] ,\w_hssi_gen3_tx_pcs_tx_test_out[7] ,\w_hssi_gen3_tx_pcs_tx_test_out[6] ,
\w_hssi_gen3_tx_pcs_tx_test_out[5] ,\w_hssi_gen3_tx_pcs_tx_test_out[4] ,\w_hssi_gen3_tx_pcs_tx_test_out[3] ,\w_hssi_gen3_tx_pcs_tx_test_out[2] ,\w_hssi_gen3_tx_pcs_tx_test_out[1] ,\w_hssi_gen3_tx_pcs_tx_test_out[0] }),
	.txdata({\w_hssi_8g_tx_pcs_tx_data_out[31] ,\w_hssi_8g_tx_pcs_tx_data_out[30] ,\w_hssi_8g_tx_pcs_tx_data_out[29] ,\w_hssi_8g_tx_pcs_tx_data_out[28] ,\w_hssi_8g_tx_pcs_tx_data_out[27] ,\w_hssi_8g_tx_pcs_tx_data_out[26] ,\w_hssi_8g_tx_pcs_tx_data_out[25] ,
\w_hssi_8g_tx_pcs_tx_data_out[24] ,\w_hssi_8g_tx_pcs_tx_data_out[23] ,\w_hssi_8g_tx_pcs_tx_data_out[22] ,\w_hssi_8g_tx_pcs_tx_data_out[21] ,\w_hssi_8g_tx_pcs_tx_data_out[20] ,\w_hssi_8g_tx_pcs_tx_data_out[19] ,\w_hssi_8g_tx_pcs_tx_data_out[18] ,
\w_hssi_8g_tx_pcs_tx_data_out[17] ,\w_hssi_8g_tx_pcs_tx_data_out[16] ,\w_hssi_8g_tx_pcs_tx_data_out[15] ,\w_hssi_8g_tx_pcs_tx_data_out[14] ,\w_hssi_8g_tx_pcs_tx_data_out[13] ,\w_hssi_8g_tx_pcs_tx_data_out[12] ,\w_hssi_8g_tx_pcs_tx_data_out[11] ,
\w_hssi_8g_tx_pcs_tx_data_out[10] ,\w_hssi_8g_tx_pcs_tx_data_out[9] ,\w_hssi_8g_tx_pcs_tx_data_out[8] ,\w_hssi_8g_tx_pcs_tx_data_out[7] ,\w_hssi_8g_tx_pcs_tx_data_out[6] ,\w_hssi_8g_tx_pcs_tx_data_out[5] ,\w_hssi_8g_tx_pcs_tx_data_out[4] ,
\w_hssi_8g_tx_pcs_tx_data_out[3] ,\w_hssi_8g_tx_pcs_tx_data_out[2] ,\w_hssi_8g_tx_pcs_tx_data_out[1] ,\w_hssi_8g_tx_pcs_tx_data_out[0] }),
	.txdatak({\w_hssi_8g_tx_pcs_tx_datak_out[3] ,\w_hssi_8g_tx_pcs_tx_datak_out[2] ,\w_hssi_8g_tx_pcs_tx_datak_out[1] ,\w_hssi_8g_tx_pcs_tx_datak_out[0] }),
	.txmargin({\w_hssi_8g_tx_pcs_phfifo_txmargin[2] ,\w_hssi_8g_tx_pcs_phfifo_txmargin[1] ,\w_hssi_8g_tx_pcs_phfifo_txmargin[0] }),
	.blockselect(out_blockselect_hssi_pipe_gen3),
	.dis_pc_byte(),
	.gen3_clk_sel(w_hssi_pipe_gen3_gen3_clk_sel),
	.pcs_rst(w_hssi_pipe_gen3_pcs_rst),
	.phystatus(w_hssi_pipe_gen3_phystatus),
	.pma_rx_det_pd(),
	.pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
	.pma_txdeemph(),
	.pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
	.pma_txswing(),
	.reset_pc_prts(),
	.rev_lpbk_8gpcs_out(w_hssi_pipe_gen3_rev_lpbk_8gpcs_out),
	.rev_lpbk_int(w_hssi_pipe_gen3_rev_lpbk_int),
	.rxelecidle(w_hssi_pipe_gen3_rxelecidle),
	.rxpolarity_8gpcs_out(w_hssi_pipe_gen3_rxpolarity_8gpcs_out),
	.rxpolarity_int(w_hssi_pipe_gen3_rxpolarity_int),
	.rxvalid(w_hssi_pipe_gen3_rxvalid),
	.shutdown_clk(w_hssi_pipe_gen3_shutdown_clk),
	.tx_blk_start_int(w_hssi_pipe_gen3_tx_blk_start_int),
	.txdataskip_int(w_hssi_pipe_gen3_txdataskip_int),
	.avmmreaddata(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_AVMMREADDATA_bus ),
	.pma_current_coeff(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_COEFF_bus ),
	.pma_current_rxpreset(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_PMA_CURRENT_RXPRESET_bus ),
	.pma_txmargin(),
	.rx_blk_start(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_BLK_START_bus ),
	.rx_sync_hdr(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RX_SYNC_HDR_bus ),
	.rxd_8gpcs_out(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXD_8GPCS_OUT_bus ),
	.rxdataskip(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXDATASKIP_bus ),
	.rxstatus(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_RXSTATUS_bus ),
	.test_out(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TEST_OUT_bus ),
	.tx_sync_hdr_int(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TX_SYNC_HDR_INT_bus ),
	.txdata_int(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATA_INT_bus ),
	.txdatak_int(\gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3_TXDATAK_INT_bus ));
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .bypass_rx_detection_enable = "false";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .bypass_rx_preset = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .bypass_rx_preset_enable = "false";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .bypass_tx_coefficent = 18'b000000000000000000;
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .bypass_tx_coefficent_enable = "false";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .elecidle_delay_g3 = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .ind_error_reporting = "dis_ind_error_reporting";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .mode = "disable_pcs";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .phy_status_delay_g12 = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .phy_status_delay_g3 = 3'b000;
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .phystatus_rst_toggle_g12 = "dis_phystatus_rst_toggle";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .phystatus_rst_toggle_g3 = "dis_phystatus_rst_toggle_g3";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .rate_match_pad_insertion = "dis_rm_fifo_pad_ins";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pipe_gen3.inst_twentynm_hssi_pipe_gen3 .test_out_sel = "disable_test_out";

twentynm_hssi_gen3_tx_pcs \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.blk_start_in(w_hssi_pipe_gen3_tx_blk_start_int),
	.data_valid(w_hssi_pipe_gen3_txdataskip_int),
	.lpbk_blk_start(w_hssi_gen3_rx_pcs_lpbk_blk_start),
	.lpbk_data_valid(w_hssi_gen3_rx_pcs_lpbk_data_valid),
	.lpbk_en(w_hssi_pipe_gen3_rev_lpbk_int),
	.tx_pma_clk(w_hssi_8g_tx_pcs_clk_out_gen3),
	.tx_rstn(w_hssi_8g_tx_pcs_g3_tx_pma_rstn),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.data_in({\w_hssi_pipe_gen3_txdata_int[31] ,\w_hssi_pipe_gen3_txdata_int[30] ,\w_hssi_pipe_gen3_txdata_int[29] ,\w_hssi_pipe_gen3_txdata_int[28] ,\w_hssi_pipe_gen3_txdata_int[27] ,\w_hssi_pipe_gen3_txdata_int[26] ,\w_hssi_pipe_gen3_txdata_int[25] ,
\w_hssi_pipe_gen3_txdata_int[24] ,\w_hssi_pipe_gen3_txdata_int[23] ,\w_hssi_pipe_gen3_txdata_int[22] ,\w_hssi_pipe_gen3_txdata_int[21] ,\w_hssi_pipe_gen3_txdata_int[20] ,\w_hssi_pipe_gen3_txdata_int[19] ,\w_hssi_pipe_gen3_txdata_int[18] ,
\w_hssi_pipe_gen3_txdata_int[17] ,\w_hssi_pipe_gen3_txdata_int[16] ,\w_hssi_pipe_gen3_txdata_int[15] ,\w_hssi_pipe_gen3_txdata_int[14] ,\w_hssi_pipe_gen3_txdata_int[13] ,\w_hssi_pipe_gen3_txdata_int[12] ,\w_hssi_pipe_gen3_txdata_int[11] ,
\w_hssi_pipe_gen3_txdata_int[10] ,\w_hssi_pipe_gen3_txdata_int[9] ,\w_hssi_pipe_gen3_txdata_int[8] ,\w_hssi_pipe_gen3_txdata_int[7] ,\w_hssi_pipe_gen3_txdata_int[6] ,\w_hssi_pipe_gen3_txdata_int[5] ,\w_hssi_pipe_gen3_txdata_int[4] ,
\w_hssi_pipe_gen3_txdata_int[3] ,\w_hssi_pipe_gen3_txdata_int[2] ,\w_hssi_pipe_gen3_txdata_int[1] ,\w_hssi_pipe_gen3_txdata_int[0] }),
	.lpbk_data_in({\w_hssi_gen3_rx_pcs_lpbk_data[33] ,\w_hssi_gen3_rx_pcs_lpbk_data[32] ,\w_hssi_gen3_rx_pcs_lpbk_data[31] ,\w_hssi_gen3_rx_pcs_lpbk_data[30] ,\w_hssi_gen3_rx_pcs_lpbk_data[29] ,\w_hssi_gen3_rx_pcs_lpbk_data[28] ,\w_hssi_gen3_rx_pcs_lpbk_data[27] ,
\w_hssi_gen3_rx_pcs_lpbk_data[26] ,\w_hssi_gen3_rx_pcs_lpbk_data[25] ,\w_hssi_gen3_rx_pcs_lpbk_data[24] ,\w_hssi_gen3_rx_pcs_lpbk_data[23] ,\w_hssi_gen3_rx_pcs_lpbk_data[22] ,\w_hssi_gen3_rx_pcs_lpbk_data[21] ,\w_hssi_gen3_rx_pcs_lpbk_data[20] ,
\w_hssi_gen3_rx_pcs_lpbk_data[19] ,\w_hssi_gen3_rx_pcs_lpbk_data[18] ,\w_hssi_gen3_rx_pcs_lpbk_data[17] ,\w_hssi_gen3_rx_pcs_lpbk_data[16] ,\w_hssi_gen3_rx_pcs_lpbk_data[15] ,\w_hssi_gen3_rx_pcs_lpbk_data[14] ,\w_hssi_gen3_rx_pcs_lpbk_data[13] ,
\w_hssi_gen3_rx_pcs_lpbk_data[12] ,\w_hssi_gen3_rx_pcs_lpbk_data[11] ,\w_hssi_gen3_rx_pcs_lpbk_data[10] ,\w_hssi_gen3_rx_pcs_lpbk_data[9] ,\w_hssi_gen3_rx_pcs_lpbk_data[8] ,\w_hssi_gen3_rx_pcs_lpbk_data[7] ,\w_hssi_gen3_rx_pcs_lpbk_data[6] ,
\w_hssi_gen3_rx_pcs_lpbk_data[5] ,\w_hssi_gen3_rx_pcs_lpbk_data[4] ,\w_hssi_gen3_rx_pcs_lpbk_data[3] ,\w_hssi_gen3_rx_pcs_lpbk_data[2] ,\w_hssi_gen3_rx_pcs_lpbk_data[1] ,\w_hssi_gen3_rx_pcs_lpbk_data[0] }),
	.sync_in({\w_hssi_pipe_gen3_tx_sync_hdr_int[1] ,\w_hssi_pipe_gen3_tx_sync_hdr_int[0] }),
	.blockselect(out_blockselect_hssi_gen3_tx_pcs),
	.avmmreaddata(\gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_AVMMREADDATA_bus ),
	.data_out(\gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_DATA_OUT_bus ),
	.par_lpbk_b4gb_out(\gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_B4GB_OUT_bus ),
	.par_lpbk_out(\gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_PAR_LPBK_OUT_bus ),
	.tx_test_out(\gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs_TX_TEST_OUT_bus ));
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .mode = "disable_pcs";
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .reverse_lpbk = "rev_lpbk_dis";
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .tx_bitslip = 5'b00000;
defparam \gen_twentynm_hssi_gen3_tx_pcs.inst_twentynm_hssi_gen3_tx_pcs .tx_gbox_byp = "bypass_gbox";

twentynm_hssi_krfec_tx_pcs \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.tx_data_valid_in(w_hssi_10g_tx_pcs_tx_data_valid_out_krfec),
	.tx_krfec_clk(w_hssi_10g_tx_pcs_tx_fec_clk),
	.tx_master_clk(w_hssi_10g_tx_pcs_tx_master_clk),
	.tx_master_clk_rst_n(w_hssi_10g_tx_pcs_tx_master_clk_rst_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.tx_control_in({\w_hssi_10g_tx_pcs_tx_control_out_krfec[8] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[7] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[6] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[5] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[4] ,
\w_hssi_10g_tx_pcs_tx_control_out_krfec[3] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[2] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[1] ,\w_hssi_10g_tx_pcs_tx_control_out_krfec[0] }),
	.tx_data_in({\w_hssi_10g_tx_pcs_tx_data_out_krfec[63] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[62] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[61] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[60] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[59] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[58] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[57] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[56] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[55] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[54] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[53] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[52] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[51] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[50] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[49] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[48] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[47] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[46] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[45] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[44] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[43] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[42] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[41] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[40] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[39] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[38] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[37] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[36] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[35] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[34] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[33] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[32] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[31] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[30] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[29] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[28] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[27] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[26] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[25] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[24] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[23] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[22] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[21] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[20] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[19] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[18] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[17] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[16] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[15] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[14] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[13] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[12] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[11] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[10] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[9] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[8] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[7] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[6] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[5] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[4] ,
\w_hssi_10g_tx_pcs_tx_data_out_krfec[3] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[2] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[1] ,\w_hssi_10g_tx_pcs_tx_data_out_krfec[0] }),
	.blockselect(out_blockselect_hssi_krfec_tx_pcs),
	.pld_10g_krfec_tx_frame_krfec_reg(),
	.pld_krfec_tx_alignment_plddirect_reg(),
	.pld_krfec_tx_alignment_reg(),
	.tx_alignment(w_hssi_krfec_tx_pcs_tx_alignment),
	.tx_frame(w_hssi_krfec_tx_pcs_tx_frame),
	.avmmreaddata(\gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_AVMMREADDATA_bus ),
	.tx_data_out(\gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_DATA_OUT_bus ),
	.tx_test_data(\gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs_TX_TEST_DATA_bus ));
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .burst_err = "burst_err_dis";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .burst_err_len = "burst_err_len1";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .ctrl_bit_reverse = "ctrl_bit_reverse_en";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .data_bit_reverse = "data_bit_reverse_dis";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .enc_frame_query = "enc_query_dis";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .low_latency_en = "disable";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .pipeln_encoder = "enable";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .pipeln_scrambler = "enable";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .prot_mode = "disable_mode";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .transcode_err = "trans_err_dis";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .transmit_order = "transmit_lsb";
defparam \gen_twentynm_hssi_krfec_tx_pcs.inst_twentynm_hssi_krfec_tx_pcs .tx_testbus_sel = "overall";

twentynm_hssi_fifo_rx_pcs \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs (
	.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.hard_reset_n(gnd),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
	.wr_clk_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_clk),
	.wr_clk_8g_clock_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_dw_clk),
	.wr_clk_8g_clock_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_rmfifo_sw_clk),
	.wr_clk_8g_phase_comp_dw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_dw_clk),
	.wr_clk_8g_phase_comp_sw(w_hssi_8g_rx_pcs_wr_clk_rx_phfifo_sw_clk),
	.wr_clk_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_clk),
	.wr_en_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_en),
	.wr_en_8g_clock_comp(w_hssi_8g_rx_pcs_wr_en_rx_rmfifo),
	.wr_en_8g_phase_comp(w_hssi_8g_rx_pcs_wr_en_rx_phfifo),
	.wr_en_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_en),
	.wr_rst_n_10g(w_hssi_10g_rx_pcs_rx_fifo_wr_rst_n),
	.wr_rst_n_8g_clock_comp(w_hssi_8g_rx_pcs_wr_rst_rx_rmfifo),
	.wr_rst_n_8g_phase_comp(w_hssi_8g_rx_pcs_wr_rst_n_rx_phfifo),
	.wr_rst_n_gen3(w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_rst_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.data_in_10g({\w_hssi_10g_rx_pcs_rx_fifo_wr_data[73] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[72] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[71] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[70] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[69] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[68] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[67] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[66] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[65] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[64] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[63] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[62] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[61] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[60] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[59] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[58] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[57] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[56] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[55] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[54] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[53] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[52] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[51] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[50] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[49] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[48] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[47] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[46] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[45] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[44] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[43] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[42] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[41] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[40] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[39] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[38] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[37] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[36] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[35] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[34] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[33] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[32] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[31] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[30] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[29] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[28] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[27] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[26] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[25] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[24] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[23] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[22] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[21] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[20] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[19] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[18] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[17] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[16] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[15] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[14] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[13] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[12] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[11] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[10] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[9] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[8] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[7] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[6] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[5] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[4] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[3] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[2] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_data[1] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_data[0] }),
	.data_in_8g_clock_comp({\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[31] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[30] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[29] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[28] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[27] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[26] ,
\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[25] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[24] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[23] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[22] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[21] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[20] ,
\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[19] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[18] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[17] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[16] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[15] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[14] ,
\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[13] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[12] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[11] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[10] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[9] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[8] ,
\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[7] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[6] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[5] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[4] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[3] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[2] ,
\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[1] ,\w_hssi_8g_rx_pcs_wr_data_rx_rmfifo[0] }),
	.data_in_8g_phase_comp({\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[79] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[78] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[77] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[76] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[75] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[74] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[73] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[72] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[71] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[70] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[69] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[68] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[67] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[66] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[65] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[64] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[63] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[62] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[61] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[60] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[59] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[58] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[57] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[56] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[55] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[54] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[53] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[52] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[51] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[50] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[49] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[48] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[47] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[46] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[45] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[44] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[43] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[42] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[41] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[40] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[39] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[38] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[37] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[36] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[35] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[34] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[33] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[32] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[31] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[30] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[29] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[28] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[27] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[26] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[25] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[24] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[23] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[22] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[21] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[20] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[19] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[18] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[17] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[16] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[15] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[14] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[13] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[12] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[11] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[10] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[9] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[8] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[7] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[6] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[5] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[4] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[3] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[2] ,
\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[1] ,\w_hssi_8g_rx_pcs_wr_data_rx_phfifo[0] }),
	.data_in_gen3({\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[39] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[38] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[37] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[36] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[35] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[34] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[33] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[32] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[31] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[30] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[29] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[28] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[27] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[26] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[25] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[24] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[23] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[22] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[21] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[20] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[19] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[18] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[17] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[16] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[15] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[14] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[13] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[12] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[11] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[10] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[9] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[8] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[7] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[6] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[5] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[4] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[3] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[2] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[1] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_data[0] }),
	.rd_ptr2_10g({\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[31] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[30] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[29] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[28] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[27] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[26] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[25] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[24] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[23] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[22] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[21] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[20] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[19] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[18] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[17] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[16] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[15] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[14] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[13] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[12] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[11] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[10] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[9] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[8] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[7] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[6] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[5] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[4] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[3] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[2] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[1] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr2[0] }),
	.rd_ptr2_8g_clock_comp({\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[19] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[18] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[17] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[16] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[15] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[14] ,
\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[13] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[12] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[11] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[10] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[9] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[8] ,
\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[7] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[6] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[5] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[4] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[3] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[2] ,
\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[1] ,\w_hssi_8g_rx_pcs_rd_ptr2_rx_rmfifo[0] }),
	.rd_ptr_10g({\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[31] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[30] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[29] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[28] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[27] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[26] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[25] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[24] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[23] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[22] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[21] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[20] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[19] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[18] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[17] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[16] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[15] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[14] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[13] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[12] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[11] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[10] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[9] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[8] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[7] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[6] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[5] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[4] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[3] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[2] ,
\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[1] ,\w_hssi_10g_rx_pcs_rx_fifo_rd_ptr[0] }),
	.rd_ptr_8g_clock_comp({\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[19] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[18] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[17] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[16] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[15] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[14] ,
\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[13] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[12] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[11] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[10] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[9] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[8] ,
\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[7] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[6] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[5] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[4] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[3] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[2] ,
\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[1] ,\w_hssi_8g_rx_pcs_rd_ptr1_rx_rmfifo[0] }),
	.rd_ptr_8g_phase_comp({\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[7] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[6] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[5] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[4] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[3] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[2] ,
\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[1] ,\w_hssi_8g_rx_pcs_rd_ptr_rx_phfifo[0] }),
	.rd_ptr_gen3({\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[15] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[14] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[13] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[12] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[11] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[10] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[9] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[8] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[7] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[6] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[5] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[4] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[3] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[2] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[1] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_rd_ptr[0] }),
	.wr_ptr_10g({\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[31] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[30] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[29] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[28] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[27] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[26] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[25] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[24] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[23] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[22] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[21] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[20] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[19] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[18] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[17] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[16] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[15] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[14] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[13] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[12] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[11] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[10] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[9] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[8] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[7] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[6] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[5] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[4] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[3] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[2] ,
\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[1] ,\w_hssi_10g_rx_pcs_rx_fifo_wr_ptr[0] }),
	.wr_ptr_8g_clock_comp({\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[19] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[18] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[17] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[16] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[15] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[14] ,
\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[13] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[12] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[11] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[10] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[9] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[8] ,
\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[7] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[6] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[5] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[4] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[3] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[2] ,
\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[1] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_rmfifo[0] }),
	.wr_ptr_8g_phase_comp({\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[7] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[6] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[5] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[4] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[3] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[2] ,
\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[1] ,\w_hssi_8g_rx_pcs_wr_ptr_rx_phfifo[0] }),
	.wr_ptr_gen3({\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[15] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[14] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[13] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[12] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[11] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[10] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[9] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[8] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[7] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[6] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[5] ,
\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[4] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[3] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[2] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[1] ,\w_hssi_gen3_rx_pcs_mem_rx_fifo_wr_ptr[0] }),
	.blockselect(out_blockselect_hssi_fifo_rx_pcs),
	.avmmreaddata(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_AVMMREADDATA_bus ),
	.data_out2_10g(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_10G_bus ),
	.data_out2_8g_clock_comp(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT2_8G_CLOCK_COMP_bus ),
	.data_out_10g(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_10G_bus ),
	.data_out_8g_clock_comp(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_CLOCK_COMP_bus ),
	.data_out_8g_phase_comp(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_8G_PHASE_COMP_bus ),
	.data_out_gen3(\gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs_DATA_OUT_GEN3_bus ));
defparam \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs .double_read_mode = "double_read_dis";
defparam \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs .prot_mode = "non_teng_mode";
defparam \gen_twentynm_hssi_fifo_rx_pcs.inst_twentynm_hssi_fifo_rx_pcs .silicon_rev = "20nm5";

twentynm_hssi_fifo_tx_pcs \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs (
	.atpg_rst_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_atpg_rst_n),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.hard_reset_n(gnd),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_mem_scan_mode_n),
	.wr_clk_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_clk),
	.wr_clk_8g_phase_comp_dw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_dw_clk),
	.wr_clk_8g_phase_comp_sw(w_hssi_8g_tx_pcs_wr_clk_tx_phfifo_sw_clk),
	.wr_en_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_en),
	.wr_en_8g_phase_comp(w_hssi_8g_tx_pcs_wr_en_tx_phfifo),
	.wr_rst_n_10g(w_hssi_10g_tx_pcs_tx_fifo_wr_rst_n),
	.wr_rst_n_8g_phase_comp(w_hssi_8g_tx_pcs_wr_rst_n_tx_phfifo),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.data_in2_10g({\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[72] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[71] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[70] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[69] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[68] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[67] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[66] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[65] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[64] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[63] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[62] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[61] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[60] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[59] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[58] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[57] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[56] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[55] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[54] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[53] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[52] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[51] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[50] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[49] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[48] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[47] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[46] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[45] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[44] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[43] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[42] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[41] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[40] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[39] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[38] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[37] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[36] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[35] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[34] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[33] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[32] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[31] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[30] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[29] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[28] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[27] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[26] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[25] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[24] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[23] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[22] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[21] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[20] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[19] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[18] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[17] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[16] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[15] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[14] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[13] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[12] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[11] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[10] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[9] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[8] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[7] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[6] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[5] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[4] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[3] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[2] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[1] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data_dw[0] }),
	.data_in_10g({\w_hssi_10g_tx_pcs_tx_fifo_wr_data[72] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[71] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[70] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[69] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[68] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[67] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[66] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[65] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[64] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[63] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[62] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[61] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[60] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[59] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[58] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[57] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[56] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[55] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[54] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[53] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[52] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[51] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[50] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[49] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[48] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[47] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[46] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[45] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[44] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[43] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[42] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[41] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[40] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[39] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[38] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[37] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[36] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[35] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[34] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[33] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[32] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[31] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[30] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[29] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[28] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[27] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[26] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[25] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[24] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[23] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[22] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[21] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[20] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[19] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[18] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[17] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[16] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[15] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[14] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[13] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[12] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[11] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[10] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[9] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[8] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[7] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[6] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[5] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[4] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[3] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[2] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_data[1] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_data[0] }),
	.data_in_8g_phase_comp({\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[63] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[62] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[61] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[60] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[59] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[58] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[57] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[56] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[55] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[54] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[53] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[52] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[51] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[50] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[49] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[48] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[47] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[46] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[45] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[44] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[43] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[42] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[41] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[40] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[39] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[38] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[37] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[36] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[35] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[34] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[33] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[32] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[31] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[30] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[29] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[28] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[27] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[26] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[25] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[24] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[23] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[22] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[21] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[20] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[19] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[18] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[17] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[16] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[15] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[14] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[13] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[12] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[11] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[10] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[9] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[8] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[7] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[6] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[5] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[4] ,
\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[3] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[2] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[1] ,\w_hssi_8g_tx_pcs_wr_data_tx_phfifo[0] }),
	.rd_ptr_10g({\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[15] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[14] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[13] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[12] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[11] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[10] ,
\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[9] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[8] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[7] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[6] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[5] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[4] ,
\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[3] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[2] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[1] ,\w_hssi_10g_tx_pcs_tx_fifo_rd_ptr[0] }),
	.rd_ptr_8g_phase_comp({\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[7] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[6] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[5] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[4] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[3] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[2] ,
\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[1] ,\w_hssi_8g_tx_pcs_rd_ptr_tx_phfifo[0] }),
	.wr_ptr_10g({\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[15] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[14] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[13] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[12] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[11] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[10] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[9] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[8] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[7] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[6] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[5] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[4] ,
\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[3] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[2] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[1] ,\w_hssi_10g_tx_pcs_tx_fifo_wr_ptr[0] }),
	.wr_ptr_8g_phase_comp({\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[7] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[6] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[5] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[4] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[3] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[2] ,
\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[1] ,\w_hssi_8g_tx_pcs_wr_ptr_tx_phfifo[0] }),
	.blockselect(out_blockselect_hssi_fifo_tx_pcs),
	.avmmreaddata(\gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_AVMMREADDATA_bus ),
	.data_out_10g(\gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_10G_bus ),
	.data_out_8g_phase_comp(\gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs_DATA_OUT_8G_PHASE_COMP_bus ));
defparam \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs .double_write_mode = "double_write_dis";
defparam \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs .prot_mode = "non_teng_mode";
defparam \gen_twentynm_hssi_fifo_tx_pcs.inst_twentynm_hssi_fifo_tx_pcs .silicon_rev = "20nm5";

twentynm_hssi_common_pcs_pma_interface \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pmaif_8g_pipe_tx_pma_rstn(w_hssi_8g_tx_pcs_pmaif_asn_rstn),
	.int_pmaif_8g_rev_lpbk(w_hssi_pipe_gen1_2_rev_loopbk),
	.int_pmaif_8g_tx_clk_out_gen3(w_hssi_8g_tx_pcs_tx_clk_out_pmaif),
	.int_pmaif_8g_txdetectrx(w_hssi_pipe_gen1_2_txdetectrx),
	.int_pmaif_g3_pma_txdetectrx(w_hssi_pipe_gen3_pma_txdetectrx),
	.int_pmaif_g3_rev_lpbk(w_hssi_pipe_gen3_rev_lpbk_int),
	.int_pmaif_pldif_8g_tx_pld_rstn(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_8g_txurstpcs_n),
	.int_pmaif_pldif_adapt_start(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_adapt_start),
	.int_pmaif_pldif_atpg_los_en_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_atpg_los_en_n),
	.int_pmaif_pldif_csr_test_dis(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_csr_test_dis),
	.int_pmaif_pldif_early_eios(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_early_eios),
	.int_pmaif_pldif_ltd_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltd_b),
	.int_pmaif_pldif_ltr(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ltr),
	.int_pmaif_pldif_nfrzdrv(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nfrzdrv),
	.int_pmaif_pldif_nrpi_freeze(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_nrpi_freeze),
	.int_pmaif_pldif_pma_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
	.int_pmaif_pldif_pma_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
	.int_pmaif_pldif_ppm_lock(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_ppm_lock),
	.int_pmaif_pldif_refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
	.int_pmaif_pldif_rs_lpbk_b(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rs_lpbk_b),
	.int_pmaif_pldif_rx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rx_qpi_pullup),
	.int_pmaif_pldif_rxpma_rstb(w_hssi_rx_pld_pcs_interface_int_pldif_pmaif_rxpma_rstb),
	.int_pmaif_pldif_tx_bitslip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bitslip),
	.int_pmaif_pldif_tx_bonding_rstb(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_bonding_rstb),
	.int_pmaif_pldif_tx_pma_syncp_hip(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_pma_syncp_hip),
	.int_pmaif_pldif_tx_qpi_pulldn(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pulldn),
	.int_pmaif_pldif_tx_qpi_pullup(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_tx_qpi_pullup),
	.int_pmaif_pldif_txdetectrx(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_txdetectrx),
	.int_pmaif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
	.int_rx_dft_obsrv_clk(w_hssi_rx_pcs_pma_interface_int_rx_dft_obsrv_clk),
	.iocsr_clk(gnd),
	.iocsr_rdy(vcc),
	.iocsr_rdy_dly(vcc),
	.pma_adapt_done(gnd),
	.pma_clklow(in_pma_clklow),
	.pma_fref(in_pma_fref),
	.pma_hclk(gnd),
	.pma_pfdmode_lock(in_pma_pfdmode_lock),
	.pma_signal_det(in_pma_signal_det),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.int_pmaif_8g_current_coeff({\w_hssi_pipe_gen1_2_current_coeff[17] ,\w_hssi_pipe_gen1_2_current_coeff[16] ,\w_hssi_pipe_gen1_2_current_coeff[15] ,\w_hssi_pipe_gen1_2_current_coeff[14] ,\w_hssi_pipe_gen1_2_current_coeff[13] ,\w_hssi_pipe_gen1_2_current_coeff[12] ,
\w_hssi_pipe_gen1_2_current_coeff[11] ,\w_hssi_pipe_gen1_2_current_coeff[10] ,\w_hssi_pipe_gen1_2_current_coeff[9] ,\w_hssi_pipe_gen1_2_current_coeff[8] ,\w_hssi_pipe_gen1_2_current_coeff[7] ,\w_hssi_pipe_gen1_2_current_coeff[6] ,
\w_hssi_pipe_gen1_2_current_coeff[5] ,\w_hssi_pipe_gen1_2_current_coeff[4] ,\w_hssi_pipe_gen1_2_current_coeff[3] ,\w_hssi_pipe_gen1_2_current_coeff[2] ,\w_hssi_pipe_gen1_2_current_coeff[1] ,\w_hssi_pipe_gen1_2_current_coeff[0] }),
	.int_pmaif_8g_eios_det({\w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[2] ,\w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[1] ,\w_hssi_8g_rx_pcs_eios_det_cdr_ctrl[0] }),
	.int_pmaif_g3_eios_det({w_hssi_gen3_rx_pcs_ei_det_int,w_hssi_gen3_rx_pcs_ei_partial_det_int,w_hssi_gen3_rx_pcs_i_det_int}),
	.int_pmaif_g3_pma_current_coeff({\w_hssi_pipe_gen3_pma_current_coeff[17] ,\w_hssi_pipe_gen3_pma_current_coeff[16] ,\w_hssi_pipe_gen3_pma_current_coeff[15] ,\w_hssi_pipe_gen3_pma_current_coeff[14] ,\w_hssi_pipe_gen3_pma_current_coeff[13] ,\w_hssi_pipe_gen3_pma_current_coeff[12] ,
\w_hssi_pipe_gen3_pma_current_coeff[11] ,\w_hssi_pipe_gen3_pma_current_coeff[10] ,\w_hssi_pipe_gen3_pma_current_coeff[9] ,\w_hssi_pipe_gen3_pma_current_coeff[8] ,\w_hssi_pipe_gen3_pma_current_coeff[7] ,\w_hssi_pipe_gen3_pma_current_coeff[6] ,
\w_hssi_pipe_gen3_pma_current_coeff[5] ,\w_hssi_pipe_gen3_pma_current_coeff[4] ,\w_hssi_pipe_gen3_pma_current_coeff[3] ,\w_hssi_pipe_gen3_pma_current_coeff[2] ,\w_hssi_pipe_gen3_pma_current_coeff[1] ,\w_hssi_pipe_gen3_pma_current_coeff[0] }),
	.int_pmaif_g3_pma_current_rxpreset({\w_hssi_pipe_gen3_pma_current_rxpreset[2] ,\w_hssi_pipe_gen3_pma_current_rxpreset[1] ,\w_hssi_pipe_gen3_pma_current_rxpreset[0] }),
	.int_pmaif_pldif_interface_select(),
	.int_pmaif_pldif_pcie_switch({\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pcie_switch[0] }),
	.int_pmaif_pldif_pma_reserved_out({\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[4] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[3] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[2] ,
\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_reserved_out[0] }),
	.int_pmaif_pldif_rate({\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[1] ,\w_hssi_common_pld_pcs_interface_int_pldif_pmaif_rate[0] }),
	.int_tx_dft_obsrv_clk({\w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[4] ,\w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[3] ,\w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[2] ,\w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[1] ,
\w_hssi_tx_pcs_pma_interface_int_tx_dft_obsrv_clk[0] }),
	.iocsr_config({gnd,gnd,gnd,gnd,gnd,gnd}),
	.pma_pcie_sw_done({in_pma_pcie_sw_done[1],in_pma_pcie_sw_done[0]}),
	.pma_reserved_in({gnd,gnd,gnd,gnd,vcc}),
	.pma_testbus({gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.pmaif_bundling_in_down({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.pmaif_bundling_in_up({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rx_pmaif_test_out({\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[19] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[18] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[17] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[16] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[15] ,
\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[14] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[13] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[12] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[11] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[10] ,
\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[9] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[8] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[7] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[6] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[5] ,
\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[4] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[3] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[2] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[1] ,\w_hssi_rx_pcs_pma_interface_rx_pmaif_test_out[0] }),
	.rx_prbs_ver_test({\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[19] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[18] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[17] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[16] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[15] ,
\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[14] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[13] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[12] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[11] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[10] ,
\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[9] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[8] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[7] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[6] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[5] ,
\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[4] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[3] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[2] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[1] ,\w_hssi_rx_pcs_pma_interface_rx_prbs_ver_test[0] }),
	.tx_prbs_gen_test({\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[19] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[18] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[17] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[16] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[15] ,
\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[14] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[13] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[12] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[11] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[10] ,
\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[9] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[8] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[7] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[6] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[5] ,
\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[4] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[3] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[2] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[1] ,\w_hssi_tx_pcs_pma_interface_tx_prbs_gen_test[0] }),
	.uhsif_test_out_1({\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[19] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[18] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[17] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[16] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[15] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[14] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[13] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[12] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[11] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[10] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[9] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[8] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[7] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[6] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[5] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[4] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[3] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[2] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[1] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_1[0] }),
	.uhsif_test_out_2({\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[19] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[18] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[17] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[16] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[15] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[14] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[13] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[12] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[11] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[10] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[9] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[8] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[7] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[6] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[5] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[4] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[3] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[2] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[1] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_2[0] }),
	.uhsif_test_out_3({\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[19] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[18] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[17] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[16] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[15] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[14] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[13] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[12] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[11] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[10] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[9] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[8] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[7] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[6] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[5] ,
\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[4] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[3] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[2] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[1] ,\w_hssi_tx_pcs_pma_interface_uhsif_test_out_3[0] }),
	.blockselect(out_blockselect_hssi_common_pcs_pma_interface),
	.int_pmaif_8g_eios_detected(w_hssi_common_pcs_pma_interface_int_pmaif_8g_eios_detected),
	.int_pmaif_8g_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_8g_inferred_rxvalid),
	.int_pmaif_8g_power_state_transition_done(w_hssi_common_pcs_pma_interface_int_pmaif_8g_power_state_transition_done),
	.int_pmaif_avmm_iocsr_clk(),
	.int_pmaif_avmm_iocsr_rdy(),
	.int_pmaif_avmm_iocsr_rdy_dly(),
	.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
	.int_pmaif_g3_inferred_rxvalid(w_hssi_common_pcs_pma_interface_int_pmaif_g3_inferred_rxvalid),
	.int_pmaif_pldif_adapt_done(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_adapt_done),
	.int_pmaif_pldif_dft_obsrv_clk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_dft_obsrv_clk),
	.int_pmaif_pldif_mask_tx_pll(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_mask_tx_pll),
	.int_pmaif_pldif_pfdmode_lock(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pfdmode_lock),
	.int_pmaif_pldif_pma_clklow(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_clklow),
	.int_pmaif_pldif_pma_fref(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_fref),
	.int_pmaif_pldif_pma_hclk(w_hssi_common_pcs_pma_interface_int_pmaif_pldif_pma_hclk),
	.pma_adapt_start(),
	.pma_atpg_los_en_n(),
	.pma_csr_test_dis(),
	.pma_early_eios(out_pma_early_eios),
	.pma_ltd_b(out_pma_ltd_b),
	.pma_ltr(out_pma_ltr),
	.pma_nfrzdrv(),
	.pma_nrpi_freeze(),
	.pma_ppm_lock(out_pma_ppm_lock),
	.pma_rs_lpbk_b(out_pma_rs_lpbk_b),
	.pma_rx_qpi_pullup(out_pma_rx_qpi_pullup),
	.pma_scan_mode_n(),
	.pma_scan_shift_n(),
	.pma_tx_bitslip(out_pma_tx_bitslip),
	.pma_tx_bonding_rstb(out_pma_tx_bonding_rstb),
	.pma_tx_pma_syncp(),
	.pma_tx_qpi_pulldn(out_pma_tx_qpi_pulldn),
	.pma_tx_qpi_pullup(out_pma_tx_qpi_pullup),
	.pma_tx_txdetectrx(out_pma_tx_txdetectrx),
	.sta_pma_hclk_by2(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface~O_STA_PMA_HCLK_BY2 ),
	.avmmreaddata(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_AVMMREADDATA_bus ),
	.int_pmaif_8g_asn_bundling_in(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_8G_ASN_BUNDLING_IN_bus ),
	.int_pmaif_avmm_iocsr_config(),
	.int_pmaif_g3_pcs_asn_bundling_in(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_G3_PCS_ASN_BUNDLING_IN_bus ),
	.int_pmaif_pldif_pcie_sw_done(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PCIE_SW_DONE_bus ),
	.int_pmaif_pldif_pma_reserved_in(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_PMA_RESERVED_IN_bus ),
	.int_pmaif_pldif_test_out(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TEST_OUT_bus ),
	.int_pmaif_pldif_testbus(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_INT_PMAIF_PLDIF_TESTBUS_bus ),
	.pma_current_coeff(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_CURRENT_COEFF_bus ),
	.pma_current_rxpreset(),
	.pma_interface_select(),
	.pma_pcie_switch(\gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface_PMA_PCIE_SWITCH_bus ),
	.pma_reserved_out(),
	.pmaif_bundling_out_down(),
	.pmaif_bundling_out_up());
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .asn_clk_enable = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .asn_enable = "dis_asn";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .block_sel = "eight_g_pcs";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_early_eios = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_pcie_switch = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_pma_ltr = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_pma_sw_done = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_ppm_lock = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_send_syncp_fbkp = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .bypass_txdetectrx = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .cdr_control = "dis_cdr_ctrl";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .cid_enable = "dis_cid_mode";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .cp_cons_sel = "cp_cons_master";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .cp_dwn_mstr = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .cp_up_mstr = "true";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ctrl_plane_bonding = "individual";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .data_mask_count = 16'b0000000000000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .data_mask_count_multi = 3'b000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .dft_observation_clock_selection = "dft_clk_obsrv_tx0";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .early_eios_counter = 8'b00000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .force_freqdet = "force_freqdet_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .free_run_clk_enable = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ignore_sigdet_g23 = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pc_en_counter = 7'b0000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pc_rst_counter = 5'b00000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pcie_hip_mode = "hip_disable";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ph_fifo_reg_mode = "phfifo_reg_mode_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .phfifo_flush_wait = 6'b000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pipe_if_g3pcs = "pipe_if_8gpcs";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pma_done_counter = 18'b000000000000000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pma_if_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .pma_if_dft_val = "dft_0";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppm_cnt_rst = "ppm_cnt_rst_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppm_deassert_early = "deassert_early_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppm_det_buckets = "ppm_100_bucket";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppm_gen1_2_cnt = "cnt_32k";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppm_post_eidle_delay = "cnt_200_cycles";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .ppmsel = "ppmsel_1000";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .prot_mode = "other_protocols";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .rxvalid_mask = "rxvalid_mask_dis";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .sigdet_wait_counter = 12'b000000000000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .sigdet_wait_counter_multi = 3'b000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .sim_mode = "disable";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .spd_chg_rst_wait_cnt_en = "false";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .testout_sel = "asn_test";
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .wait_clk_on_off_timer = 4'b0000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .wait_pipe_synchronizing = 5'b00000;
defparam \gen_twentynm_hssi_common_pcs_pma_interface.inst_twentynm_hssi_common_pcs_pma_interface .wait_send_syncp_fbkp = 11'b00000000000;

twentynm_hssi_tx_pcs_pma_interface \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.int_pmaif_10g_tx_clk_out(w_hssi_10g_tx_pcs_tx_clk_out_pma_if),
	.int_pmaif_8g_tx_clk_out(w_hssi_8g_tx_pcs_tx_clk_out_8g_pmaif),
	.int_pmaif_8g_tx_elec_idle(w_hssi_pipe_gen1_2_tx_elec_idle_out),
	.int_pmaif_g3_data_sel(w_hssi_common_pcs_pma_interface_int_pmaif_g3_data_sel),
	.int_pmaif_g3_pma_tx_elec_idle(w_hssi_pipe_gen3_pma_tx_elec_idle),
	.int_pmaif_pldif_pmaif_tx_pld_rst_n(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_pld_rst_n),
	.int_pmaif_pldif_polinv_tx(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_polinv_tx),
	.int_pmaif_pldif_txelecidle(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txelecidle),
	.int_pmaif_pldif_txpma_rstb(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_txpma_rstb),
	.int_pmaif_pldif_uhsif_scan_chain_in(w_hssi_common_pld_pcs_interface_int_pmaif_pldif_uhsif_scan_chain_in),
	.int_pmaif_pldif_uhsif_tx_clk(w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_clk),
	.pma_tx_clkdiv_user(in_pma_tx_clkdiv_user),
	.pma_tx_pma_clk(in_pma_tx_pma_clk),
	.refclk_dig(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_refclk_dig),
	.refclk_dig_uhsif(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_uhsif_refclk_dig),
	.scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_scan_mode_n),
	.uhsif_scan_mode_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_mode_n),
	.uhsif_scan_shift_n(w_hssi_common_pld_pcs_interface_int_pldif_pmaif_pma_scan_shift_n),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.int_pmaif_10g_tx_pma_data({\w_hssi_10g_tx_pcs_tx_pma_data[63] ,\w_hssi_10g_tx_pcs_tx_pma_data[62] ,\w_hssi_10g_tx_pcs_tx_pma_data[61] ,\w_hssi_10g_tx_pcs_tx_pma_data[60] ,\w_hssi_10g_tx_pcs_tx_pma_data[59] ,\w_hssi_10g_tx_pcs_tx_pma_data[58] ,\w_hssi_10g_tx_pcs_tx_pma_data[57] ,
\w_hssi_10g_tx_pcs_tx_pma_data[56] ,\w_hssi_10g_tx_pcs_tx_pma_data[55] ,\w_hssi_10g_tx_pcs_tx_pma_data[54] ,\w_hssi_10g_tx_pcs_tx_pma_data[53] ,\w_hssi_10g_tx_pcs_tx_pma_data[52] ,\w_hssi_10g_tx_pcs_tx_pma_data[51] ,\w_hssi_10g_tx_pcs_tx_pma_data[50] ,
\w_hssi_10g_tx_pcs_tx_pma_data[49] ,\w_hssi_10g_tx_pcs_tx_pma_data[48] ,\w_hssi_10g_tx_pcs_tx_pma_data[47] ,\w_hssi_10g_tx_pcs_tx_pma_data[46] ,\w_hssi_10g_tx_pcs_tx_pma_data[45] ,\w_hssi_10g_tx_pcs_tx_pma_data[44] ,\w_hssi_10g_tx_pcs_tx_pma_data[43] ,
\w_hssi_10g_tx_pcs_tx_pma_data[42] ,\w_hssi_10g_tx_pcs_tx_pma_data[41] ,\w_hssi_10g_tx_pcs_tx_pma_data[40] ,\w_hssi_10g_tx_pcs_tx_pma_data[39] ,\w_hssi_10g_tx_pcs_tx_pma_data[38] ,\w_hssi_10g_tx_pcs_tx_pma_data[37] ,\w_hssi_10g_tx_pcs_tx_pma_data[36] ,
\w_hssi_10g_tx_pcs_tx_pma_data[35] ,\w_hssi_10g_tx_pcs_tx_pma_data[34] ,\w_hssi_10g_tx_pcs_tx_pma_data[33] ,\w_hssi_10g_tx_pcs_tx_pma_data[32] ,\w_hssi_10g_tx_pcs_tx_pma_data[31] ,\w_hssi_10g_tx_pcs_tx_pma_data[30] ,\w_hssi_10g_tx_pcs_tx_pma_data[29] ,
\w_hssi_10g_tx_pcs_tx_pma_data[28] ,\w_hssi_10g_tx_pcs_tx_pma_data[27] ,\w_hssi_10g_tx_pcs_tx_pma_data[26] ,\w_hssi_10g_tx_pcs_tx_pma_data[25] ,\w_hssi_10g_tx_pcs_tx_pma_data[24] ,\w_hssi_10g_tx_pcs_tx_pma_data[23] ,\w_hssi_10g_tx_pcs_tx_pma_data[22] ,
\w_hssi_10g_tx_pcs_tx_pma_data[21] ,\w_hssi_10g_tx_pcs_tx_pma_data[20] ,\w_hssi_10g_tx_pcs_tx_pma_data[19] ,\w_hssi_10g_tx_pcs_tx_pma_data[18] ,\w_hssi_10g_tx_pcs_tx_pma_data[17] ,\w_hssi_10g_tx_pcs_tx_pma_data[16] ,\w_hssi_10g_tx_pcs_tx_pma_data[15] ,
\w_hssi_10g_tx_pcs_tx_pma_data[14] ,\w_hssi_10g_tx_pcs_tx_pma_data[13] ,\w_hssi_10g_tx_pcs_tx_pma_data[12] ,\w_hssi_10g_tx_pcs_tx_pma_data[11] ,\w_hssi_10g_tx_pcs_tx_pma_data[10] ,\w_hssi_10g_tx_pcs_tx_pma_data[9] ,\w_hssi_10g_tx_pcs_tx_pma_data[8] ,
\w_hssi_10g_tx_pcs_tx_pma_data[7] ,\w_hssi_10g_tx_pcs_tx_pma_data[6] ,\w_hssi_10g_tx_pcs_tx_pma_data[5] ,\w_hssi_10g_tx_pcs_tx_pma_data[4] ,\w_hssi_10g_tx_pcs_tx_pma_data[3] ,\w_hssi_10g_tx_pcs_tx_pma_data[2] ,\w_hssi_10g_tx_pcs_tx_pma_data[1] ,
\w_hssi_10g_tx_pcs_tx_pma_data[0] }),
	.int_pmaif_10g_tx_pma_data_gate_val({\w_hssi_10g_tx_pcs_tx_pma_gating_val[63] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[62] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[61] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[60] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[59] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[58] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[57] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[56] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[55] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[54] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[53] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[52] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[51] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[50] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[49] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[48] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[47] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[46] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[45] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[44] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[43] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[42] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[41] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[40] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[39] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[38] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[37] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[36] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[35] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[34] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[33] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[32] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[31] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[30] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[29] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[28] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[27] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[26] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[25] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[24] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[23] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[22] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[21] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[20] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[19] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[18] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[17] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[16] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[15] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[14] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[13] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[12] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[11] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[10] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[9] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[8] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[7] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[6] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[5] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[4] ,
\w_hssi_10g_tx_pcs_tx_pma_gating_val[3] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[2] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[1] ,\w_hssi_10g_tx_pcs_tx_pma_gating_val[0] }),
	.int_pmaif_8g_pudr({\w_hssi_8g_tx_pcs_dataout[19] ,\w_hssi_8g_tx_pcs_dataout[18] ,\w_hssi_8g_tx_pcs_dataout[17] ,\w_hssi_8g_tx_pcs_dataout[16] ,\w_hssi_8g_tx_pcs_dataout[15] ,\w_hssi_8g_tx_pcs_dataout[14] ,\w_hssi_8g_tx_pcs_dataout[13] ,\w_hssi_8g_tx_pcs_dataout[12] ,
\w_hssi_8g_tx_pcs_dataout[11] ,\w_hssi_8g_tx_pcs_dataout[10] ,\w_hssi_8g_tx_pcs_dataout[9] ,\w_hssi_8g_tx_pcs_dataout[8] ,\w_hssi_8g_tx_pcs_dataout[7] ,\w_hssi_8g_tx_pcs_dataout[6] ,\w_hssi_8g_tx_pcs_dataout[5] ,\w_hssi_8g_tx_pcs_dataout[4] ,
\w_hssi_8g_tx_pcs_dataout[3] ,\w_hssi_8g_tx_pcs_dataout[2] ,\w_hssi_8g_tx_pcs_dataout[1] ,\w_hssi_8g_tx_pcs_dataout[0] }),
	.int_pmaif_g3_pma_data_out({\w_hssi_gen3_tx_pcs_data_out[31] ,\w_hssi_gen3_tx_pcs_data_out[30] ,\w_hssi_gen3_tx_pcs_data_out[29] ,\w_hssi_gen3_tx_pcs_data_out[28] ,\w_hssi_gen3_tx_pcs_data_out[27] ,\w_hssi_gen3_tx_pcs_data_out[26] ,\w_hssi_gen3_tx_pcs_data_out[25] ,
\w_hssi_gen3_tx_pcs_data_out[24] ,\w_hssi_gen3_tx_pcs_data_out[23] ,\w_hssi_gen3_tx_pcs_data_out[22] ,\w_hssi_gen3_tx_pcs_data_out[21] ,\w_hssi_gen3_tx_pcs_data_out[20] ,\w_hssi_gen3_tx_pcs_data_out[19] ,\w_hssi_gen3_tx_pcs_data_out[18] ,
\w_hssi_gen3_tx_pcs_data_out[17] ,\w_hssi_gen3_tx_pcs_data_out[16] ,\w_hssi_gen3_tx_pcs_data_out[15] ,\w_hssi_gen3_tx_pcs_data_out[14] ,\w_hssi_gen3_tx_pcs_data_out[13] ,\w_hssi_gen3_tx_pcs_data_out[12] ,\w_hssi_gen3_tx_pcs_data_out[11] ,
\w_hssi_gen3_tx_pcs_data_out[10] ,\w_hssi_gen3_tx_pcs_data_out[9] ,\w_hssi_gen3_tx_pcs_data_out[8] ,\w_hssi_gen3_tx_pcs_data_out[7] ,\w_hssi_gen3_tx_pcs_data_out[6] ,\w_hssi_gen3_tx_pcs_data_out[5] ,\w_hssi_gen3_tx_pcs_data_out[4] ,
\w_hssi_gen3_tx_pcs_data_out[3] ,\w_hssi_gen3_tx_pcs_data_out[2] ,\w_hssi_gen3_tx_pcs_data_out[1] ,\w_hssi_gen3_tx_pcs_data_out[0] }),
	.int_pmaif_pldif_tx_data({\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[63] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[62] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[61] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[60] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[59] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[58] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[57] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[56] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[55] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[54] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[53] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[52] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[51] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[50] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[49] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[48] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[47] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[46] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[45] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[44] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[40] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[39] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[36] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[34] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[32] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[29] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[28] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[20] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[19] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[16] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[14] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[12] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[8] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_tx_data[0] }),
	.int_pmaif_pldif_uhsif_tx_data({\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[63] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[62] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[61] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[60] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[59] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[58] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[57] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[56] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[55] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[54] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[53] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[52] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[51] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[50] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[49] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[48] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[47] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[46] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[45] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[44] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[43] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[42] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[41] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[40] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[39] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[38] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[37] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[36] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[35] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[34] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[33] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[32] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[31] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[30] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[29] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[28] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[27] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[26] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[25] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[24] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[23] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[22] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[21] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[20] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[19] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[18] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[17] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[16] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[15] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[14] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[13] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[12] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[11] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[10] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[9] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[8] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[7] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[6] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[5] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[4] ,
\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[3] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[2] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[1] ,\w_hssi_tx_pld_pcs_interface_int_pldif_pmaif_uhsif_tx_data[0] }),
	.write_en(),
	.blockselect(out_blockselect_hssi_tx_pcs_pma_interface),
	.int_pmaif_10g_tx_pma_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_10g_tx_pma_clk),
	.int_pmaif_8g_txpma_local_clk(w_hssi_tx_pcs_pma_interface_int_pmaif_8g_txpma_local_clk),
	.int_pmaif_pldif_tx_clkdiv(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv),
	.int_pmaif_pldif_tx_clkdiv_user(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_tx_clkdiv_user),
	.int_pmaif_pldif_uhsif_lock(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_lock),
	.int_pmaif_pldif_uhsif_scan_chain_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_scan_chain_out),
	.int_pmaif_pldif_uhsif_tx_clk_out(w_hssi_tx_pcs_pma_interface_int_pmaif_pldif_uhsif_tx_clk_out),
	.pma_tx_elec_idle(out_pma_tx_elec_idle),
	.pma_txpma_rstb(out_pma_txpma_rstb),
	.avmm_user_dataout(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMM_USER_DATAOUT_bus ),
	.avmmreaddata(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_AVMMREADDATA_bus ),
	.int_tx_dft_obsrv_clk(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_INT_TX_DFT_OBSRV_CLK_bus ),
	.pma_tx_pma_data(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_PMA_TX_PMA_DATA_bus ),
	.tx_pma_data_loopback(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_DATA_LOOPBACK_bus ),
	.tx_pma_uhsif_data_loopback(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PMA_UHSIF_DATA_LOOPBACK_bus ),
	.tx_prbs_gen_test(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_TX_PRBS_GEN_TEST_bus ),
	.uhsif_test_out_1(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_1_bus ),
	.uhsif_test_out_2(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_2_bus ),
	.uhsif_test_out_3(\gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface_UHSIF_TEST_OUT_3_bus ),
	.write_en_ack());
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .bypass_pma_txelecidle = "true";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .channel_operation_mode = "tx_rx_pair_enabled";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .lpbk_en = "disable";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .master_clk_sel = "master_tx_pma_clk";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .pcie_sub_prot_mode_tx = "other_prot_mode";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .pldif_datawidth_mode = "pldif_data_10bit";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .pma_dw_tx = "pma_10b_tx";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .pma_if_dft_en = "dft_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .pmagate_en = "pmagate_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .prbs9_dwidth = "prbs9_64b";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .prbs_clken = "prbs_clk_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .prbs_gen_pat = "prbs_gen_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .prot_mode_tx = "eightg_only_pld_mode_tx";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .reconfig_settings = "{}";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .sq_wave_num = "sq_wave_default";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .sqwgen_clken = "sqwgen_clk_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .tx_dyn_polarity_inversion = "tx_dyn_polinv_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .tx_pma_data_sel = "eight_g_pcs";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .tx_static_polarity_inversion = "tx_stat_polinv_dis";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_cnt_step_filt_before_lock = "uhsif_filt_stepsz_b4lock_2";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_cnt_thresh_filt_after_lock_value = 4'b0000;
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_cnt_thresh_filt_before_lock = "uhsif_filt_cntthr_b4lock_8";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dcn_test_update_period = "uhsif_dcn_test_period_4";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dcn_testmode_enable = "uhsif_dcn_test_mode_disable";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dead_zone_count_thresh = "uhsif_dzt_cnt_thr_2";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dead_zone_detection_enable = "uhsif_dzt_disable";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dead_zone_obser_window = "uhsif_dzt_obr_win_16";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dead_zone_skip_size = "uhsif_dzt_skipsz_4";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_delay_cell_index_sel = "uhsif_index_cram";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_delay_cell_margin = "uhsif_dcn_margin_2";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_delay_cell_static_index_value = 8'b00000000;
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dft_dead_zone_control = "uhsif_dft_dz_det_val_0";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_dft_up_filt_control = "uhsif_dft_up_val_0";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_enable = "uhsif_disable";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_segsz_after_lock = "uhsif_lkd_segsz_aflock_512";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_segsz_before_lock = "uhsif_lkd_segsz_b4lock_16";
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_thresh_cnt_after_lock_value = 4'b0000;
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_thresh_cnt_before_lock_value = 4'b0000;
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_thresh_diff_after_lock_value = 4'b0000;
defparam \gen_twentynm_hssi_tx_pcs_pma_interface.inst_twentynm_hssi_tx_pcs_pma_interface .uhsif_lock_det_thresh_diff_before_lock_value = 4'b0000;

endmodule

module wr_arria10_e3p1_det_phy_twentynm_pma_rev_20nm5 (
	in_avmmclk,
	in_avmmread,
	in_avmmrstn,
	in_avmmwrite,
	in_avmmaddress,
	in_avmmwritedata,
	out_blockselect_pma_tx_buf,
	out_rx_detect_valid,
	out_rx_found,
	out_tx_p,
	out_avmmreaddata_pma_tx_buf,
	in_rx_bitslip,
	in_rx_pma_rstb,
	in_eye_monitor,
	out_blockselect_pma_tx_ser,
	out_iqtxrxclk_out1,
	out_clkdiv_tx_user,
	out_avmmreaddata_pma_tx_ser,
	out_blockselect_pma_cgb,
	out_avmmreaddata_pma_cgb,
	out_pcie_sw_done,
	out_blockselect_pma_rx_deser,
	out_clkdiv_rx,
	out_clkdiv_rx_user,
	out_avmmreaddata_pma_rx_deser,
	out_rxdata,
	out_blockselect_pma_rx_buf,
	out_avmmreaddata_pma_rx_buf,
	out_blockselect_pma_rx_sd,
	out_sd,
	out_avmmreaddata_pma_rx_sd,
	out_blockselect_pma_rx_odi,
	out_avmmreaddata_pma_rx_odi,
	out_blockselect_pma_rx_dfe,
	out_avmmreaddata_pma_rx_dfe,
	out_blockselect_cdr_pll,
	out_clklow,
	out_fref,
	out_pfdmode_lock,
	out_rxpll_lock,
	out_avmmreaddata_cdr_pll,
	out_blockselect_pma_cdr_refclk,
	out_avmmreaddata_pma_cdr_refclk,
	out_blockselect_pma_adapt,
	out_avmmreaddata_pma_adapt,
	in_early_eios,
	in_ltd_b,
	in_ltr,
	in_ppm_lock,
	in_rs_lpbk_b,
	in_rx_qpi_pulldn,
	in_tx_bitslip,
	in_tx_bonding_rstb,
	in_tx_qpi_pulldn,
	in_tx_qpi_pullup,
	in_tx_det_rx,
	in_i_coeff,
	in_pcie_sw,
	in_tx_elec_idle,
	in_tx_pma_rstb,
	in_tx_data,
	in_rx_p,
	in_clk_fpll_b,
	in_ref_iqclk)/* synthesis synthesis_greybox=1 */;
input 	in_avmmclk;
input 	in_avmmread;
input 	in_avmmrstn;
input 	in_avmmwrite;
input 	[8:0] in_avmmaddress;
input 	[7:0] in_avmmwritedata;
output 	out_blockselect_pma_tx_buf;
output 	out_rx_detect_valid;
output 	out_rx_found;
output 	out_tx_p;
output 	[7:0] out_avmmreaddata_pma_tx_buf;
input 	in_rx_bitslip;
input 	in_rx_pma_rstb;
input 	[5:0] in_eye_monitor;
output 	out_blockselect_pma_tx_ser;
output 	out_iqtxrxclk_out1;
output 	out_clkdiv_tx_user;
output 	[7:0] out_avmmreaddata_pma_tx_ser;
output 	out_blockselect_pma_cgb;
output 	[7:0] out_avmmreaddata_pma_cgb;
output 	[1:0] out_pcie_sw_done;
output 	out_blockselect_pma_rx_deser;
output 	out_clkdiv_rx;
output 	out_clkdiv_rx_user;
output 	[7:0] out_avmmreaddata_pma_rx_deser;
output 	[63:0] out_rxdata;
output 	out_blockselect_pma_rx_buf;
output 	[7:0] out_avmmreaddata_pma_rx_buf;
output 	out_blockselect_pma_rx_sd;
output 	out_sd;
output 	[7:0] out_avmmreaddata_pma_rx_sd;
output 	out_blockselect_pma_rx_odi;
output 	[7:0] out_avmmreaddata_pma_rx_odi;
output 	out_blockselect_pma_rx_dfe;
output 	[7:0] out_avmmreaddata_pma_rx_dfe;
output 	out_blockselect_cdr_pll;
output 	out_clklow;
output 	out_fref;
output 	out_pfdmode_lock;
output 	out_rxpll_lock;
output 	[7:0] out_avmmreaddata_cdr_pll;
output 	out_blockselect_pma_cdr_refclk;
output 	[7:0] out_avmmreaddata_pma_cdr_refclk;
output 	out_blockselect_pma_adapt;
output 	[7:0] out_avmmreaddata_pma_adapt;
input 	in_early_eios;
input 	in_ltd_b;
input 	in_ltr;
input 	in_ppm_lock;
input 	in_rs_lpbk_b;
input 	in_rx_qpi_pulldn;
input 	in_tx_bitslip;
input 	in_tx_bonding_rstb;
input 	in_tx_qpi_pulldn;
input 	in_tx_qpi_pullup;
input 	in_tx_det_rx;
input 	[17:0] in_i_coeff;
input 	[1:0] in_pcie_sw;
input 	in_tx_elec_idle;
input 	in_tx_pma_rstb;
input 	[63:0] in_tx_data;
input 	in_rx_p;
input 	in_clk_fpll_b;
input 	[11:0] in_ref_iqclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \w_pma_tx_buf_atbsel[0] ;
wire \w_pma_tx_buf_atbsel[1] ;
wire \w_pma_tx_buf_atbsel[2] ;
wire \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi~atb0 ;
wire \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll~O_CDR_LPBKDP ;
wire w_pma_tx_buf_ckn;
wire w_pma_tx_buf_ckp;
wire w_pma_tx_buf_lbvon;
wire w_pma_tx_buf_lbvop;
wire w_pma_tx_ser_ckdrvn;
wire w_pma_tx_ser_ckdrvp;
wire w_pma_tx_ser_oe;
wire w_pma_tx_ser_oeb;
wire w_pma_tx_ser_oo;
wire w_pma_tx_ser_oob;
wire w_pma_cgb_bitslipstate;
wire w_pma_cgb_div2;
wire w_pma_cgb_div4;
wire w_pma_cgb_div5;
wire w_pma_cgb_hifreqclkn;
wire w_pma_cgb_hifreqclkp;
wire w_pma_cgb_rstb;
wire \w_pma_cgb_cpulse_out_bus[0] ;
wire \w_pma_cgb_cpulse_out_bus[1] ;
wire \w_pma_cgb_cpulse_out_bus[2] ;
wire \w_pma_cgb_cpulse_out_bus[3] ;
wire \w_pma_cgb_cpulse_out_bus[4] ;
wire \w_pma_cgb_cpulse_out_bus[5] ;
wire \w_pma_cgb_pcie_sw_master[1] ;
wire w_pma_rx_deser_adapt_clk;
wire w_pma_rx_deser_clkdivrx_rx;
wire \w_pma_rx_deser_data[0] ;
wire \w_pma_rx_deser_data[1] ;
wire \w_pma_rx_deser_data[2] ;
wire \w_pma_rx_deser_data[3] ;
wire \w_pma_rx_deser_data[4] ;
wire \w_pma_rx_deser_data[5] ;
wire \w_pma_rx_deser_data[6] ;
wire \w_pma_rx_deser_data[7] ;
wire \w_pma_rx_deser_data[8] ;
wire \w_pma_rx_deser_data[9] ;
wire \w_pma_rx_deser_data[10] ;
wire \w_pma_rx_deser_data[11] ;
wire \w_pma_rx_deser_data[12] ;
wire \w_pma_rx_deser_data[13] ;
wire \w_pma_rx_deser_data[14] ;
wire \w_pma_rx_deser_data[15] ;
wire \w_pma_rx_deser_data[16] ;
wire \w_pma_rx_deser_data[17] ;
wire \w_pma_rx_deser_data[18] ;
wire \w_pma_rx_deser_data[19] ;
wire \w_pma_rx_deser_data[20] ;
wire \w_pma_rx_deser_data[21] ;
wire \w_pma_rx_deser_data[22] ;
wire \w_pma_rx_deser_data[23] ;
wire \w_pma_rx_deser_data[24] ;
wire \w_pma_rx_deser_data[25] ;
wire \w_pma_rx_deser_data[26] ;
wire \w_pma_rx_deser_data[27] ;
wire \w_pma_rx_deser_data[28] ;
wire \w_pma_rx_deser_data[29] ;
wire \w_pma_rx_deser_data[30] ;
wire \w_pma_rx_deser_data[31] ;
wire \w_pma_rx_deser_data[32] ;
wire \w_pma_rx_deser_data[33] ;
wire \w_pma_rx_deser_data[34] ;
wire \w_pma_rx_deser_data[35] ;
wire \w_pma_rx_deser_data[36] ;
wire \w_pma_rx_deser_data[37] ;
wire \w_pma_rx_deser_data[38] ;
wire \w_pma_rx_deser_data[39] ;
wire \w_pma_rx_deser_data[40] ;
wire \w_pma_rx_deser_data[41] ;
wire \w_pma_rx_deser_data[42] ;
wire \w_pma_rx_deser_data[43] ;
wire \w_pma_rx_deser_data[44] ;
wire \w_pma_rx_deser_data[45] ;
wire \w_pma_rx_deser_data[46] ;
wire \w_pma_rx_deser_data[47] ;
wire \w_pma_rx_deser_data[48] ;
wire \w_pma_rx_deser_data[49] ;
wire \w_pma_rx_deser_data[50] ;
wire \w_pma_rx_deser_data[51] ;
wire \w_pma_rx_deser_data[52] ;
wire \w_pma_rx_deser_data[53] ;
wire \w_pma_rx_deser_data[54] ;
wire \w_pma_rx_deser_data[55] ;
wire \w_pma_rx_deser_data[56] ;
wire \w_pma_rx_deser_data[57] ;
wire \w_pma_rx_deser_data[58] ;
wire \w_pma_rx_deser_data[59] ;
wire \w_pma_rx_deser_data[60] ;
wire \w_pma_rx_deser_data[61] ;
wire \w_pma_rx_deser_data[62] ;
wire \w_pma_rx_deser_data[63] ;
wire \w_pma_rx_deser_error_deser[0] ;
wire \w_pma_rx_deser_error_deser[1] ;
wire \w_pma_rx_deser_error_deser[2] ;
wire \w_pma_rx_deser_error_deser[3] ;
wire \w_pma_rx_deser_error_deser[4] ;
wire \w_pma_rx_deser_error_deser[5] ;
wire \w_pma_rx_deser_error_deser[6] ;
wire \w_pma_rx_deser_error_deser[7] ;
wire \w_pma_rx_deser_error_deser[8] ;
wire \w_pma_rx_deser_error_deser[9] ;
wire \w_pma_rx_deser_error_deser[10] ;
wire \w_pma_rx_deser_error_deser[11] ;
wire \w_pma_rx_deser_error_deser[12] ;
wire \w_pma_rx_deser_error_deser[13] ;
wire \w_pma_rx_deser_error_deser[14] ;
wire \w_pma_rx_deser_error_deser[15] ;
wire \w_pma_rx_deser_error_deser[16] ;
wire \w_pma_rx_deser_error_deser[17] ;
wire \w_pma_rx_deser_error_deser[18] ;
wire \w_pma_rx_deser_error_deser[19] ;
wire \w_pma_rx_deser_error_deser[20] ;
wire \w_pma_rx_deser_error_deser[21] ;
wire \w_pma_rx_deser_error_deser[22] ;
wire \w_pma_rx_deser_error_deser[23] ;
wire \w_pma_rx_deser_error_deser[24] ;
wire \w_pma_rx_deser_error_deser[25] ;
wire \w_pma_rx_deser_error_deser[26] ;
wire \w_pma_rx_deser_error_deser[27] ;
wire \w_pma_rx_deser_error_deser[28] ;
wire \w_pma_rx_deser_error_deser[29] ;
wire \w_pma_rx_deser_error_deser[30] ;
wire \w_pma_rx_deser_error_deser[31] ;
wire \w_pma_rx_deser_error_deser[32] ;
wire \w_pma_rx_deser_error_deser[33] ;
wire \w_pma_rx_deser_error_deser[34] ;
wire \w_pma_rx_deser_error_deser[35] ;
wire \w_pma_rx_deser_error_deser[36] ;
wire \w_pma_rx_deser_error_deser[37] ;
wire \w_pma_rx_deser_error_deser[38] ;
wire \w_pma_rx_deser_error_deser[39] ;
wire \w_pma_rx_deser_error_deser[40] ;
wire \w_pma_rx_deser_error_deser[41] ;
wire \w_pma_rx_deser_error_deser[42] ;
wire \w_pma_rx_deser_error_deser[43] ;
wire \w_pma_rx_deser_error_deser[44] ;
wire \w_pma_rx_deser_error_deser[45] ;
wire \w_pma_rx_deser_error_deser[46] ;
wire \w_pma_rx_deser_error_deser[47] ;
wire \w_pma_rx_deser_error_deser[48] ;
wire \w_pma_rx_deser_error_deser[49] ;
wire \w_pma_rx_deser_error_deser[50] ;
wire \w_pma_rx_deser_error_deser[51] ;
wire \w_pma_rx_deser_error_deser[52] ;
wire \w_pma_rx_deser_error_deser[53] ;
wire \w_pma_rx_deser_error_deser[54] ;
wire \w_pma_rx_deser_error_deser[55] ;
wire \w_pma_rx_deser_error_deser[56] ;
wire \w_pma_rx_deser_error_deser[57] ;
wire \w_pma_rx_deser_error_deser[58] ;
wire \w_pma_rx_deser_error_deser[59] ;
wire \w_pma_rx_deser_error_deser[60] ;
wire \w_pma_rx_deser_error_deser[61] ;
wire \w_pma_rx_deser_error_deser[62] ;
wire \w_pma_rx_deser_error_deser[63] ;
wire \w_pma_rx_deser_odi_dout[0] ;
wire \w_pma_rx_deser_odi_dout[1] ;
wire \w_pma_rx_deser_odi_dout[2] ;
wire \w_pma_rx_deser_odi_dout[3] ;
wire \w_pma_rx_deser_odi_dout[4] ;
wire \w_pma_rx_deser_odi_dout[5] ;
wire \w_pma_rx_deser_odi_dout[6] ;
wire \w_pma_rx_deser_odi_dout[7] ;
wire \w_pma_rx_deser_odi_dout[8] ;
wire \w_pma_rx_deser_odi_dout[9] ;
wire \w_pma_rx_deser_odi_dout[10] ;
wire \w_pma_rx_deser_odi_dout[11] ;
wire \w_pma_rx_deser_odi_dout[12] ;
wire \w_pma_rx_deser_odi_dout[13] ;
wire \w_pma_rx_deser_odi_dout[14] ;
wire \w_pma_rx_deser_odi_dout[15] ;
wire \w_pma_rx_deser_odi_dout[16] ;
wire \w_pma_rx_deser_odi_dout[17] ;
wire \w_pma_rx_deser_odi_dout[18] ;
wire \w_pma_rx_deser_odi_dout[19] ;
wire \w_pma_rx_deser_odi_dout[20] ;
wire \w_pma_rx_deser_odi_dout[21] ;
wire \w_pma_rx_deser_odi_dout[22] ;
wire \w_pma_rx_deser_odi_dout[23] ;
wire \w_pma_rx_deser_odi_dout[24] ;
wire \w_pma_rx_deser_odi_dout[25] ;
wire \w_pma_rx_deser_odi_dout[26] ;
wire \w_pma_rx_deser_odi_dout[27] ;
wire \w_pma_rx_deser_odi_dout[28] ;
wire \w_pma_rx_deser_odi_dout[29] ;
wire \w_pma_rx_deser_odi_dout[30] ;
wire \w_pma_rx_deser_odi_dout[31] ;
wire \w_pma_rx_deser_odi_dout[32] ;
wire \w_pma_rx_deser_odi_dout[33] ;
wire \w_pma_rx_deser_odi_dout[34] ;
wire \w_pma_rx_deser_odi_dout[35] ;
wire \w_pma_rx_deser_odi_dout[36] ;
wire \w_pma_rx_deser_odi_dout[37] ;
wire \w_pma_rx_deser_odi_dout[38] ;
wire \w_pma_rx_deser_odi_dout[39] ;
wire \w_pma_rx_deser_odi_dout[40] ;
wire \w_pma_rx_deser_odi_dout[41] ;
wire \w_pma_rx_deser_odi_dout[42] ;
wire \w_pma_rx_deser_odi_dout[43] ;
wire \w_pma_rx_deser_odi_dout[44] ;
wire \w_pma_rx_deser_odi_dout[45] ;
wire \w_pma_rx_deser_odi_dout[46] ;
wire \w_pma_rx_deser_odi_dout[47] ;
wire \w_pma_rx_deser_odi_dout[48] ;
wire \w_pma_rx_deser_odi_dout[49] ;
wire \w_pma_rx_deser_odi_dout[50] ;
wire \w_pma_rx_deser_odi_dout[51] ;
wire \w_pma_rx_deser_odi_dout[52] ;
wire \w_pma_rx_deser_odi_dout[53] ;
wire \w_pma_rx_deser_odi_dout[54] ;
wire \w_pma_rx_deser_odi_dout[55] ;
wire \w_pma_rx_deser_odi_dout[56] ;
wire \w_pma_rx_deser_odi_dout[57] ;
wire \w_pma_rx_deser_odi_dout[58] ;
wire \w_pma_rx_deser_odi_dout[59] ;
wire \w_pma_rx_deser_odi_dout[60] ;
wire \w_pma_rx_deser_odi_dout[61] ;
wire \w_pma_rx_deser_odi_dout[62] ;
wire \w_pma_rx_deser_odi_dout[63] ;
wire \w_pma_rx_deser_pcie_sw_ret[0] ;
wire \w_pma_rx_deser_pcie_sw_ret[1] ;
wire w_pma_rx_buf_inn;
wire w_pma_rx_buf_inp;
wire w_pma_rx_buf_outn;
wire w_pma_rx_buf_outp;
wire w_pma_rx_buf_pull_dn;
wire w_pma_rx_buf_rdlpbkn;
wire w_pma_rx_buf_rdlpbkp;
wire w_pma_rx_odi_clk0_eye;
wire w_pma_rx_odi_clk0_eye_lb;
wire w_pma_rx_odi_clk180_eye;
wire w_pma_rx_odi_clk180_eye_lb;
wire w_pma_rx_odi_de_eye;
wire w_pma_rx_odi_deb_eye;
wire w_pma_rx_odi_do_eye;
wire w_pma_rx_odi_dob_eye;
wire w_pma_rx_odi_odi_en;
wire w_pma_rx_dfe_clk0_bbpd;
wire w_pma_rx_dfe_clk180_bbpd;
wire w_pma_rx_dfe_clk270_bbpd;
wire w_pma_rx_dfe_clk90_bbpd;
wire w_pma_rx_dfe_deven;
wire w_pma_rx_dfe_devenb;
wire w_pma_rx_dfe_dodd;
wire w_pma_rx_dfe_doddb;
wire w_pma_rx_dfe_edge270;
wire w_pma_rx_dfe_edge270b;
wire w_pma_rx_dfe_edge90;
wire w_pma_rx_dfe_edge90b;
wire w_pma_rx_dfe_err_ev;
wire w_pma_rx_dfe_err_evb;
wire w_pma_rx_dfe_err_od;
wire w_pma_rx_dfe_err_odb;
wire w_pma_rx_dfe_spec_vrefh;
wire w_pma_rx_dfe_spec_vrefl;
wire w_cdr_pll_clk0_des;
wire w_cdr_pll_clk0_odi;
wire w_cdr_pll_clk0_pd;
wire w_cdr_pll_clk0_pfd;
wire w_cdr_pll_clk180_des;
wire w_cdr_pll_clk180_odi;
wire w_cdr_pll_clk180_pd;
wire w_cdr_pll_clk180_pfd;
wire w_cdr_pll_clk270_odi;
wire w_cdr_pll_clk270_pd;
wire w_cdr_pll_clk90_odi;
wire w_cdr_pll_clk90_pd;
wire w_cdr_pll_deven_des;
wire w_cdr_pll_devenb_des;
wire w_cdr_pll_dodd_des;
wire w_cdr_pll_doddb_des;
wire w_cdr_pll_error_even_des;
wire w_cdr_pll_error_evenb_des;
wire w_cdr_pll_error_odd_des;
wire w_cdr_pll_error_oddb_des;
wire w_cdr_pll_rlpbkdn;
wire w_cdr_pll_rlpbkdp;
wire w_cdr_pll_rlpbkn;
wire w_cdr_pll_rlpbkp;
wire w_cdr_pll_tx_rlpbk;
wire w_pma_cdr_refclk_refclk;
wire w_pma_cdr_refclk_rx_det_clk;
wire w_pma_adapt_dfe_adapt_en;
wire w_pma_adapt_dfe_adp_clk;
wire w_pma_adapt_dfe_fltap1_sgn;
wire w_pma_adapt_dfe_fltap2_sgn;
wire w_pma_adapt_dfe_fltap3_sgn;
wire w_pma_adapt_dfe_fltap4_sgn;
wire w_pma_adapt_dfe_fltap_bypdeser;
wire w_pma_adapt_dfe_fxtap2_sgn;
wire w_pma_adapt_dfe_fxtap3_sgn;
wire w_pma_adapt_dfe_fxtap4_sgn;
wire w_pma_adapt_dfe_fxtap5_sgn;
wire w_pma_adapt_dfe_fxtap6_sgn;
wire w_pma_adapt_dfe_fxtap7_sgn;
wire w_pma_adapt_dfe_spec_disable;
wire w_pma_adapt_dfe_spec_sign_sel;
wire w_pma_adapt_dfe_vref_sign_sel;
wire \w_pma_adapt_ctle_acgain_4s[0] ;
wire \w_pma_adapt_ctle_acgain_4s[1] ;
wire \w_pma_adapt_ctle_acgain_4s[2] ;
wire \w_pma_adapt_ctle_acgain_4s[3] ;
wire \w_pma_adapt_ctle_acgain_4s[4] ;
wire \w_pma_adapt_ctle_acgain_4s[5] ;
wire \w_pma_adapt_ctle_acgain_4s[6] ;
wire \w_pma_adapt_ctle_acgain_4s[7] ;
wire \w_pma_adapt_ctle_acgain_4s[8] ;
wire \w_pma_adapt_ctle_acgain_4s[9] ;
wire \w_pma_adapt_ctle_acgain_4s[10] ;
wire \w_pma_adapt_ctle_acgain_4s[11] ;
wire \w_pma_adapt_ctle_acgain_4s[12] ;
wire \w_pma_adapt_ctle_acgain_4s[13] ;
wire \w_pma_adapt_ctle_acgain_4s[14] ;
wire \w_pma_adapt_ctle_acgain_4s[15] ;
wire \w_pma_adapt_ctle_acgain_4s[16] ;
wire \w_pma_adapt_ctle_acgain_4s[17] ;
wire \w_pma_adapt_ctle_acgain_4s[18] ;
wire \w_pma_adapt_ctle_acgain_4s[19] ;
wire \w_pma_adapt_ctle_acgain_4s[20] ;
wire \w_pma_adapt_ctle_acgain_4s[21] ;
wire \w_pma_adapt_ctle_acgain_4s[22] ;
wire \w_pma_adapt_ctle_acgain_4s[23] ;
wire \w_pma_adapt_ctle_acgain_4s[24] ;
wire \w_pma_adapt_ctle_acgain_4s[25] ;
wire \w_pma_adapt_ctle_acgain_4s[26] ;
wire \w_pma_adapt_ctle_acgain_4s[27] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[0] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[1] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[2] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[3] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[4] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[5] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[6] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[7] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[8] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[9] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[10] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[11] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[12] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[13] ;
wire \w_pma_adapt_ctle_eqz_1s_sel[14] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[0] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[1] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[2] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[3] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[4] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[5] ;
wire \w_pma_adapt_ctle_lfeq_fb_sel[6] ;
wire \w_pma_adapt_dfe_fltap1[0] ;
wire \w_pma_adapt_dfe_fltap1[1] ;
wire \w_pma_adapt_dfe_fltap1[2] ;
wire \w_pma_adapt_dfe_fltap1[3] ;
wire \w_pma_adapt_dfe_fltap1[4] ;
wire \w_pma_adapt_dfe_fltap1[5] ;
wire \w_pma_adapt_dfe_fltap2[0] ;
wire \w_pma_adapt_dfe_fltap2[1] ;
wire \w_pma_adapt_dfe_fltap2[2] ;
wire \w_pma_adapt_dfe_fltap2[3] ;
wire \w_pma_adapt_dfe_fltap2[4] ;
wire \w_pma_adapt_dfe_fltap2[5] ;
wire \w_pma_adapt_dfe_fltap3[0] ;
wire \w_pma_adapt_dfe_fltap3[1] ;
wire \w_pma_adapt_dfe_fltap3[2] ;
wire \w_pma_adapt_dfe_fltap3[3] ;
wire \w_pma_adapt_dfe_fltap3[4] ;
wire \w_pma_adapt_dfe_fltap3[5] ;
wire \w_pma_adapt_dfe_fltap4[0] ;
wire \w_pma_adapt_dfe_fltap4[1] ;
wire \w_pma_adapt_dfe_fltap4[2] ;
wire \w_pma_adapt_dfe_fltap4[3] ;
wire \w_pma_adapt_dfe_fltap4[4] ;
wire \w_pma_adapt_dfe_fltap4[5] ;
wire \w_pma_adapt_dfe_fltap_position[0] ;
wire \w_pma_adapt_dfe_fltap_position[1] ;
wire \w_pma_adapt_dfe_fltap_position[2] ;
wire \w_pma_adapt_dfe_fltap_position[3] ;
wire \w_pma_adapt_dfe_fltap_position[4] ;
wire \w_pma_adapt_dfe_fltap_position[5] ;
wire \w_pma_adapt_dfe_fxtap1[0] ;
wire \w_pma_adapt_dfe_fxtap1[1] ;
wire \w_pma_adapt_dfe_fxtap1[2] ;
wire \w_pma_adapt_dfe_fxtap1[3] ;
wire \w_pma_adapt_dfe_fxtap1[4] ;
wire \w_pma_adapt_dfe_fxtap1[5] ;
wire \w_pma_adapt_dfe_fxtap1[6] ;
wire \w_pma_adapt_dfe_fxtap2[0] ;
wire \w_pma_adapt_dfe_fxtap2[1] ;
wire \w_pma_adapt_dfe_fxtap2[2] ;
wire \w_pma_adapt_dfe_fxtap2[3] ;
wire \w_pma_adapt_dfe_fxtap2[4] ;
wire \w_pma_adapt_dfe_fxtap2[5] ;
wire \w_pma_adapt_dfe_fxtap2[6] ;
wire \w_pma_adapt_dfe_fxtap3[0] ;
wire \w_pma_adapt_dfe_fxtap3[1] ;
wire \w_pma_adapt_dfe_fxtap3[2] ;
wire \w_pma_adapt_dfe_fxtap3[3] ;
wire \w_pma_adapt_dfe_fxtap3[4] ;
wire \w_pma_adapt_dfe_fxtap3[5] ;
wire \w_pma_adapt_dfe_fxtap3[6] ;
wire \w_pma_adapt_dfe_fxtap4[0] ;
wire \w_pma_adapt_dfe_fxtap4[1] ;
wire \w_pma_adapt_dfe_fxtap4[2] ;
wire \w_pma_adapt_dfe_fxtap4[3] ;
wire \w_pma_adapt_dfe_fxtap4[4] ;
wire \w_pma_adapt_dfe_fxtap4[5] ;
wire \w_pma_adapt_dfe_fxtap5[0] ;
wire \w_pma_adapt_dfe_fxtap5[1] ;
wire \w_pma_adapt_dfe_fxtap5[2] ;
wire \w_pma_adapt_dfe_fxtap5[3] ;
wire \w_pma_adapt_dfe_fxtap5[4] ;
wire \w_pma_adapt_dfe_fxtap5[5] ;
wire \w_pma_adapt_dfe_fxtap6[0] ;
wire \w_pma_adapt_dfe_fxtap6[1] ;
wire \w_pma_adapt_dfe_fxtap6[2] ;
wire \w_pma_adapt_dfe_fxtap6[3] ;
wire \w_pma_adapt_dfe_fxtap6[4] ;
wire \w_pma_adapt_dfe_fxtap7[0] ;
wire \w_pma_adapt_dfe_fxtap7[1] ;
wire \w_pma_adapt_dfe_fxtap7[2] ;
wire \w_pma_adapt_dfe_fxtap7[3] ;
wire \w_pma_adapt_dfe_fxtap7[4] ;
wire \w_pma_adapt_odi_vref[0] ;
wire \w_pma_adapt_odi_vref[1] ;
wire \w_pma_adapt_odi_vref[2] ;
wire \w_pma_adapt_odi_vref[3] ;
wire \w_pma_adapt_odi_vref[4] ;
wire \w_pma_adapt_vga_sel[0] ;
wire \w_pma_adapt_vga_sel[1] ;
wire \w_pma_adapt_vga_sel[2] ;
wire \w_pma_adapt_vga_sel[3] ;
wire \w_pma_adapt_vga_sel[4] ;
wire \w_pma_adapt_vga_sel[5] ;
wire \w_pma_adapt_vga_sel[6] ;
wire \w_pma_adapt_vref_sel[0] ;
wire \w_pma_adapt_vref_sel[1] ;
wire \w_pma_adapt_vref_sel[2] ;
wire \w_pma_adapt_vref_sel[3] ;
wire \w_pma_adapt_vref_sel[4] ;

wire [7:0] \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus ;
wire [2:0] \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_ATBSEL_bus ;
wire [7:0] \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus ;
wire [5:0] \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus ;
wire [1:0] \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_DONE_bus ;
wire [1:0] \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_MASTER_bus ;
wire [63:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus ;
wire [7:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus ;
wire [63:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus ;
wire [63:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus ;
wire [63:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus ;
wire [1:0] \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_PCIE_SW_RET_bus ;
wire [7:0] \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus ;
wire [7:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus ;
wire [27:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus ;
wire [14:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus ;
wire [6:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus ;
wire [6:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus ;
wire [6:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus ;
wire [6:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus ;
wire [5:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus ;
wire [4:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus ;
wire [4:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus ;
wire [4:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus ;
wire [6:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus ;
wire [4:0] \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus ;

assign out_avmmreaddata_pma_tx_buf[0] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_tx_buf[1] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_tx_buf[2] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_tx_buf[3] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_tx_buf[4] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_tx_buf[5] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_tx_buf[6] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_tx_buf[7] = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus [7];

assign \w_pma_tx_buf_atbsel[0]  = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_ATBSEL_bus [0];
assign \w_pma_tx_buf_atbsel[1]  = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_ATBSEL_bus [1];
assign \w_pma_tx_buf_atbsel[2]  = \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_ATBSEL_bus [2];

assign out_avmmreaddata_pma_tx_ser[0] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_tx_ser[1] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_tx_ser[2] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_tx_ser[3] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_tx_ser[4] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_tx_ser[5] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_tx_ser[6] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_tx_ser[7] = \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_cgb[0] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_cgb[1] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_cgb[2] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_cgb[3] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_cgb[4] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_cgb[5] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_cgb[6] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_cgb[7] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus [7];

assign \w_pma_cgb_cpulse_out_bus[0]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [0];
assign \w_pma_cgb_cpulse_out_bus[1]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [1];
assign \w_pma_cgb_cpulse_out_bus[2]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [2];
assign \w_pma_cgb_cpulse_out_bus[3]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [3];
assign \w_pma_cgb_cpulse_out_bus[4]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [4];
assign \w_pma_cgb_cpulse_out_bus[5]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus [5];

assign out_pcie_sw_done[0] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_DONE_bus [0];
assign out_pcie_sw_done[1] = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_DONE_bus [1];

assign \w_pma_cgb_pcie_sw_master[1]  = \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_MASTER_bus [1];

assign out_rxdata[0] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [0];
assign out_rxdata[1] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [1];
assign out_rxdata[2] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [2];
assign out_rxdata[3] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [3];
assign out_rxdata[4] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [4];
assign out_rxdata[5] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [5];
assign out_rxdata[6] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [6];
assign out_rxdata[7] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [7];
assign out_rxdata[8] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [8];
assign out_rxdata[9] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [9];
assign out_rxdata[10] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [10];
assign out_rxdata[11] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [11];
assign out_rxdata[12] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [12];
assign out_rxdata[13] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [13];
assign out_rxdata[14] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [14];
assign out_rxdata[15] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [15];
assign out_rxdata[16] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [16];
assign out_rxdata[17] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [17];
assign out_rxdata[18] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [18];
assign out_rxdata[19] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [19];
assign out_rxdata[20] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [20];
assign out_rxdata[21] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [21];
assign out_rxdata[22] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [22];
assign out_rxdata[23] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [23];
assign out_rxdata[24] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [24];
assign out_rxdata[25] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [25];
assign out_rxdata[26] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [26];
assign out_rxdata[27] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [27];
assign out_rxdata[28] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [28];
assign out_rxdata[29] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [29];
assign out_rxdata[30] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [30];
assign out_rxdata[31] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [31];
assign out_rxdata[32] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [32];
assign out_rxdata[33] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [33];
assign out_rxdata[34] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [34];
assign out_rxdata[35] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [35];
assign out_rxdata[36] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [36];
assign out_rxdata[37] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [37];
assign out_rxdata[38] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [38];
assign out_rxdata[39] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [39];
assign out_rxdata[40] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [40];
assign out_rxdata[41] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [41];
assign out_rxdata[42] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [42];
assign out_rxdata[43] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [43];
assign out_rxdata[44] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [44];
assign out_rxdata[45] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [45];
assign out_rxdata[46] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [46];
assign out_rxdata[47] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [47];
assign out_rxdata[48] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [48];
assign out_rxdata[49] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [49];
assign out_rxdata[50] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [50];
assign out_rxdata[51] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [51];
assign out_rxdata[52] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [52];
assign out_rxdata[53] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [53];
assign out_rxdata[54] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [54];
assign out_rxdata[55] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [55];
assign out_rxdata[56] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [56];
assign out_rxdata[57] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [57];
assign out_rxdata[58] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [58];
assign out_rxdata[59] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [59];
assign out_rxdata[60] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [60];
assign out_rxdata[61] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [61];
assign out_rxdata[62] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [62];
assign out_rxdata[63] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus [63];

assign out_avmmreaddata_pma_rx_deser[0] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_rx_deser[1] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_rx_deser[2] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_rx_deser[3] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_rx_deser[4] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_rx_deser[5] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_rx_deser[6] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_rx_deser[7] = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus [7];

assign \w_pma_rx_deser_data[0]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [0];
assign \w_pma_rx_deser_data[1]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [1];
assign \w_pma_rx_deser_data[2]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [2];
assign \w_pma_rx_deser_data[3]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [3];
assign \w_pma_rx_deser_data[4]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [4];
assign \w_pma_rx_deser_data[5]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [5];
assign \w_pma_rx_deser_data[6]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [6];
assign \w_pma_rx_deser_data[7]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [7];
assign \w_pma_rx_deser_data[8]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [8];
assign \w_pma_rx_deser_data[9]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [9];
assign \w_pma_rx_deser_data[10]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [10];
assign \w_pma_rx_deser_data[11]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [11];
assign \w_pma_rx_deser_data[12]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [12];
assign \w_pma_rx_deser_data[13]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [13];
assign \w_pma_rx_deser_data[14]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [14];
assign \w_pma_rx_deser_data[15]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [15];
assign \w_pma_rx_deser_data[16]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [16];
assign \w_pma_rx_deser_data[17]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [17];
assign \w_pma_rx_deser_data[18]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [18];
assign \w_pma_rx_deser_data[19]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [19];
assign \w_pma_rx_deser_data[20]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [20];
assign \w_pma_rx_deser_data[21]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [21];
assign \w_pma_rx_deser_data[22]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [22];
assign \w_pma_rx_deser_data[23]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [23];
assign \w_pma_rx_deser_data[24]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [24];
assign \w_pma_rx_deser_data[25]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [25];
assign \w_pma_rx_deser_data[26]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [26];
assign \w_pma_rx_deser_data[27]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [27];
assign \w_pma_rx_deser_data[28]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [28];
assign \w_pma_rx_deser_data[29]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [29];
assign \w_pma_rx_deser_data[30]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [30];
assign \w_pma_rx_deser_data[31]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [31];
assign \w_pma_rx_deser_data[32]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [32];
assign \w_pma_rx_deser_data[33]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [33];
assign \w_pma_rx_deser_data[34]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [34];
assign \w_pma_rx_deser_data[35]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [35];
assign \w_pma_rx_deser_data[36]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [36];
assign \w_pma_rx_deser_data[37]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [37];
assign \w_pma_rx_deser_data[38]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [38];
assign \w_pma_rx_deser_data[39]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [39];
assign \w_pma_rx_deser_data[40]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [40];
assign \w_pma_rx_deser_data[41]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [41];
assign \w_pma_rx_deser_data[42]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [42];
assign \w_pma_rx_deser_data[43]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [43];
assign \w_pma_rx_deser_data[44]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [44];
assign \w_pma_rx_deser_data[45]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [45];
assign \w_pma_rx_deser_data[46]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [46];
assign \w_pma_rx_deser_data[47]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [47];
assign \w_pma_rx_deser_data[48]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [48];
assign \w_pma_rx_deser_data[49]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [49];
assign \w_pma_rx_deser_data[50]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [50];
assign \w_pma_rx_deser_data[51]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [51];
assign \w_pma_rx_deser_data[52]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [52];
assign \w_pma_rx_deser_data[53]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [53];
assign \w_pma_rx_deser_data[54]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [54];
assign \w_pma_rx_deser_data[55]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [55];
assign \w_pma_rx_deser_data[56]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [56];
assign \w_pma_rx_deser_data[57]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [57];
assign \w_pma_rx_deser_data[58]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [58];
assign \w_pma_rx_deser_data[59]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [59];
assign \w_pma_rx_deser_data[60]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [60];
assign \w_pma_rx_deser_data[61]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [61];
assign \w_pma_rx_deser_data[62]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [62];
assign \w_pma_rx_deser_data[63]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus [63];

assign \w_pma_rx_deser_error_deser[0]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [0];
assign \w_pma_rx_deser_error_deser[1]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [1];
assign \w_pma_rx_deser_error_deser[2]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [2];
assign \w_pma_rx_deser_error_deser[3]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [3];
assign \w_pma_rx_deser_error_deser[4]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [4];
assign \w_pma_rx_deser_error_deser[5]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [5];
assign \w_pma_rx_deser_error_deser[6]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [6];
assign \w_pma_rx_deser_error_deser[7]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [7];
assign \w_pma_rx_deser_error_deser[8]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [8];
assign \w_pma_rx_deser_error_deser[9]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [9];
assign \w_pma_rx_deser_error_deser[10]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [10];
assign \w_pma_rx_deser_error_deser[11]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [11];
assign \w_pma_rx_deser_error_deser[12]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [12];
assign \w_pma_rx_deser_error_deser[13]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [13];
assign \w_pma_rx_deser_error_deser[14]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [14];
assign \w_pma_rx_deser_error_deser[15]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [15];
assign \w_pma_rx_deser_error_deser[16]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [16];
assign \w_pma_rx_deser_error_deser[17]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [17];
assign \w_pma_rx_deser_error_deser[18]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [18];
assign \w_pma_rx_deser_error_deser[19]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [19];
assign \w_pma_rx_deser_error_deser[20]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [20];
assign \w_pma_rx_deser_error_deser[21]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [21];
assign \w_pma_rx_deser_error_deser[22]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [22];
assign \w_pma_rx_deser_error_deser[23]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [23];
assign \w_pma_rx_deser_error_deser[24]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [24];
assign \w_pma_rx_deser_error_deser[25]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [25];
assign \w_pma_rx_deser_error_deser[26]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [26];
assign \w_pma_rx_deser_error_deser[27]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [27];
assign \w_pma_rx_deser_error_deser[28]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [28];
assign \w_pma_rx_deser_error_deser[29]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [29];
assign \w_pma_rx_deser_error_deser[30]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [30];
assign \w_pma_rx_deser_error_deser[31]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [31];
assign \w_pma_rx_deser_error_deser[32]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [32];
assign \w_pma_rx_deser_error_deser[33]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [33];
assign \w_pma_rx_deser_error_deser[34]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [34];
assign \w_pma_rx_deser_error_deser[35]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [35];
assign \w_pma_rx_deser_error_deser[36]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [36];
assign \w_pma_rx_deser_error_deser[37]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [37];
assign \w_pma_rx_deser_error_deser[38]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [38];
assign \w_pma_rx_deser_error_deser[39]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [39];
assign \w_pma_rx_deser_error_deser[40]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [40];
assign \w_pma_rx_deser_error_deser[41]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [41];
assign \w_pma_rx_deser_error_deser[42]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [42];
assign \w_pma_rx_deser_error_deser[43]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [43];
assign \w_pma_rx_deser_error_deser[44]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [44];
assign \w_pma_rx_deser_error_deser[45]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [45];
assign \w_pma_rx_deser_error_deser[46]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [46];
assign \w_pma_rx_deser_error_deser[47]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [47];
assign \w_pma_rx_deser_error_deser[48]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [48];
assign \w_pma_rx_deser_error_deser[49]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [49];
assign \w_pma_rx_deser_error_deser[50]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [50];
assign \w_pma_rx_deser_error_deser[51]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [51];
assign \w_pma_rx_deser_error_deser[52]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [52];
assign \w_pma_rx_deser_error_deser[53]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [53];
assign \w_pma_rx_deser_error_deser[54]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [54];
assign \w_pma_rx_deser_error_deser[55]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [55];
assign \w_pma_rx_deser_error_deser[56]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [56];
assign \w_pma_rx_deser_error_deser[57]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [57];
assign \w_pma_rx_deser_error_deser[58]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [58];
assign \w_pma_rx_deser_error_deser[59]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [59];
assign \w_pma_rx_deser_error_deser[60]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [60];
assign \w_pma_rx_deser_error_deser[61]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [61];
assign \w_pma_rx_deser_error_deser[62]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [62];
assign \w_pma_rx_deser_error_deser[63]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus [63];

assign \w_pma_rx_deser_odi_dout[0]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [0];
assign \w_pma_rx_deser_odi_dout[1]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [1];
assign \w_pma_rx_deser_odi_dout[2]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [2];
assign \w_pma_rx_deser_odi_dout[3]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [3];
assign \w_pma_rx_deser_odi_dout[4]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [4];
assign \w_pma_rx_deser_odi_dout[5]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [5];
assign \w_pma_rx_deser_odi_dout[6]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [6];
assign \w_pma_rx_deser_odi_dout[7]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [7];
assign \w_pma_rx_deser_odi_dout[8]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [8];
assign \w_pma_rx_deser_odi_dout[9]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [9];
assign \w_pma_rx_deser_odi_dout[10]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [10];
assign \w_pma_rx_deser_odi_dout[11]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [11];
assign \w_pma_rx_deser_odi_dout[12]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [12];
assign \w_pma_rx_deser_odi_dout[13]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [13];
assign \w_pma_rx_deser_odi_dout[14]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [14];
assign \w_pma_rx_deser_odi_dout[15]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [15];
assign \w_pma_rx_deser_odi_dout[16]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [16];
assign \w_pma_rx_deser_odi_dout[17]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [17];
assign \w_pma_rx_deser_odi_dout[18]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [18];
assign \w_pma_rx_deser_odi_dout[19]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [19];
assign \w_pma_rx_deser_odi_dout[20]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [20];
assign \w_pma_rx_deser_odi_dout[21]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [21];
assign \w_pma_rx_deser_odi_dout[22]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [22];
assign \w_pma_rx_deser_odi_dout[23]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [23];
assign \w_pma_rx_deser_odi_dout[24]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [24];
assign \w_pma_rx_deser_odi_dout[25]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [25];
assign \w_pma_rx_deser_odi_dout[26]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [26];
assign \w_pma_rx_deser_odi_dout[27]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [27];
assign \w_pma_rx_deser_odi_dout[28]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [28];
assign \w_pma_rx_deser_odi_dout[29]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [29];
assign \w_pma_rx_deser_odi_dout[30]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [30];
assign \w_pma_rx_deser_odi_dout[31]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [31];
assign \w_pma_rx_deser_odi_dout[32]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [32];
assign \w_pma_rx_deser_odi_dout[33]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [33];
assign \w_pma_rx_deser_odi_dout[34]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [34];
assign \w_pma_rx_deser_odi_dout[35]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [35];
assign \w_pma_rx_deser_odi_dout[36]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [36];
assign \w_pma_rx_deser_odi_dout[37]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [37];
assign \w_pma_rx_deser_odi_dout[38]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [38];
assign \w_pma_rx_deser_odi_dout[39]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [39];
assign \w_pma_rx_deser_odi_dout[40]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [40];
assign \w_pma_rx_deser_odi_dout[41]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [41];
assign \w_pma_rx_deser_odi_dout[42]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [42];
assign \w_pma_rx_deser_odi_dout[43]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [43];
assign \w_pma_rx_deser_odi_dout[44]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [44];
assign \w_pma_rx_deser_odi_dout[45]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [45];
assign \w_pma_rx_deser_odi_dout[46]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [46];
assign \w_pma_rx_deser_odi_dout[47]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [47];
assign \w_pma_rx_deser_odi_dout[48]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [48];
assign \w_pma_rx_deser_odi_dout[49]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [49];
assign \w_pma_rx_deser_odi_dout[50]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [50];
assign \w_pma_rx_deser_odi_dout[51]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [51];
assign \w_pma_rx_deser_odi_dout[52]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [52];
assign \w_pma_rx_deser_odi_dout[53]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [53];
assign \w_pma_rx_deser_odi_dout[54]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [54];
assign \w_pma_rx_deser_odi_dout[55]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [55];
assign \w_pma_rx_deser_odi_dout[56]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [56];
assign \w_pma_rx_deser_odi_dout[57]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [57];
assign \w_pma_rx_deser_odi_dout[58]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [58];
assign \w_pma_rx_deser_odi_dout[59]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [59];
assign \w_pma_rx_deser_odi_dout[60]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [60];
assign \w_pma_rx_deser_odi_dout[61]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [61];
assign \w_pma_rx_deser_odi_dout[62]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [62];
assign \w_pma_rx_deser_odi_dout[63]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus [63];

assign \w_pma_rx_deser_pcie_sw_ret[0]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_PCIE_SW_RET_bus [0];
assign \w_pma_rx_deser_pcie_sw_ret[1]  = \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_PCIE_SW_RET_bus [1];

assign out_avmmreaddata_pma_rx_buf[0] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_rx_buf[1] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_rx_buf[2] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_rx_buf[3] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_rx_buf[4] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_rx_buf[5] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_rx_buf[6] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_rx_buf[7] = \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_rx_sd[0] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_rx_sd[1] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_rx_sd[2] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_rx_sd[3] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_rx_sd[4] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_rx_sd[5] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_rx_sd[6] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_rx_sd[7] = \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_rx_odi[0] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_rx_odi[1] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_rx_odi[2] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_rx_odi[3] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_rx_odi[4] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_rx_odi[5] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_rx_odi[6] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_rx_odi[7] = \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_rx_dfe[0] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_rx_dfe[1] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_rx_dfe[2] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_rx_dfe[3] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_rx_dfe[4] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_rx_dfe[5] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_rx_dfe[6] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_rx_dfe[7] = \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus [7];

assign out_avmmreaddata_cdr_pll[0] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [0];
assign out_avmmreaddata_cdr_pll[1] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [1];
assign out_avmmreaddata_cdr_pll[2] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [2];
assign out_avmmreaddata_cdr_pll[3] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [3];
assign out_avmmreaddata_cdr_pll[4] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [4];
assign out_avmmreaddata_cdr_pll[5] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [5];
assign out_avmmreaddata_cdr_pll[6] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [6];
assign out_avmmreaddata_cdr_pll[7] = \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_cdr_refclk[0] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_cdr_refclk[1] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_cdr_refclk[2] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_cdr_refclk[3] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_cdr_refclk[4] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_cdr_refclk[5] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_cdr_refclk[6] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_cdr_refclk[7] = \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus [7];

assign out_avmmreaddata_pma_adapt[0] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [0];
assign out_avmmreaddata_pma_adapt[1] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [1];
assign out_avmmreaddata_pma_adapt[2] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [2];
assign out_avmmreaddata_pma_adapt[3] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [3];
assign out_avmmreaddata_pma_adapt[4] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [4];
assign out_avmmreaddata_pma_adapt[5] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [5];
assign out_avmmreaddata_pma_adapt[6] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [6];
assign out_avmmreaddata_pma_adapt[7] = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus [7];

assign \w_pma_adapt_ctle_acgain_4s[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [0];
assign \w_pma_adapt_ctle_acgain_4s[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [1];
assign \w_pma_adapt_ctle_acgain_4s[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [2];
assign \w_pma_adapt_ctle_acgain_4s[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [3];
assign \w_pma_adapt_ctle_acgain_4s[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [4];
assign \w_pma_adapt_ctle_acgain_4s[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [5];
assign \w_pma_adapt_ctle_acgain_4s[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [6];
assign \w_pma_adapt_ctle_acgain_4s[7]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [7];
assign \w_pma_adapt_ctle_acgain_4s[8]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [8];
assign \w_pma_adapt_ctle_acgain_4s[9]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [9];
assign \w_pma_adapt_ctle_acgain_4s[10]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [10];
assign \w_pma_adapt_ctle_acgain_4s[11]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [11];
assign \w_pma_adapt_ctle_acgain_4s[12]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [12];
assign \w_pma_adapt_ctle_acgain_4s[13]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [13];
assign \w_pma_adapt_ctle_acgain_4s[14]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [14];
assign \w_pma_adapt_ctle_acgain_4s[15]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [15];
assign \w_pma_adapt_ctle_acgain_4s[16]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [16];
assign \w_pma_adapt_ctle_acgain_4s[17]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [17];
assign \w_pma_adapt_ctle_acgain_4s[18]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [18];
assign \w_pma_adapt_ctle_acgain_4s[19]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [19];
assign \w_pma_adapt_ctle_acgain_4s[20]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [20];
assign \w_pma_adapt_ctle_acgain_4s[21]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [21];
assign \w_pma_adapt_ctle_acgain_4s[22]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [22];
assign \w_pma_adapt_ctle_acgain_4s[23]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [23];
assign \w_pma_adapt_ctle_acgain_4s[24]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [24];
assign \w_pma_adapt_ctle_acgain_4s[25]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [25];
assign \w_pma_adapt_ctle_acgain_4s[26]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [26];
assign \w_pma_adapt_ctle_acgain_4s[27]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus [27];

assign \w_pma_adapt_ctle_eqz_1s_sel[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [0];
assign \w_pma_adapt_ctle_eqz_1s_sel[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [1];
assign \w_pma_adapt_ctle_eqz_1s_sel[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [2];
assign \w_pma_adapt_ctle_eqz_1s_sel[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [3];
assign \w_pma_adapt_ctle_eqz_1s_sel[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [4];
assign \w_pma_adapt_ctle_eqz_1s_sel[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [5];
assign \w_pma_adapt_ctle_eqz_1s_sel[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [6];
assign \w_pma_adapt_ctle_eqz_1s_sel[7]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [7];
assign \w_pma_adapt_ctle_eqz_1s_sel[8]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [8];
assign \w_pma_adapt_ctle_eqz_1s_sel[9]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [9];
assign \w_pma_adapt_ctle_eqz_1s_sel[10]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [10];
assign \w_pma_adapt_ctle_eqz_1s_sel[11]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [11];
assign \w_pma_adapt_ctle_eqz_1s_sel[12]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [12];
assign \w_pma_adapt_ctle_eqz_1s_sel[13]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [13];
assign \w_pma_adapt_ctle_eqz_1s_sel[14]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus [14];

assign \w_pma_adapt_ctle_lfeq_fb_sel[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [0];
assign \w_pma_adapt_ctle_lfeq_fb_sel[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [1];
assign \w_pma_adapt_ctle_lfeq_fb_sel[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [2];
assign \w_pma_adapt_ctle_lfeq_fb_sel[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [3];
assign \w_pma_adapt_ctle_lfeq_fb_sel[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [4];
assign \w_pma_adapt_ctle_lfeq_fb_sel[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [5];
assign \w_pma_adapt_ctle_lfeq_fb_sel[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus [6];

assign \w_pma_adapt_dfe_fltap1[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [0];
assign \w_pma_adapt_dfe_fltap1[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [1];
assign \w_pma_adapt_dfe_fltap1[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [2];
assign \w_pma_adapt_dfe_fltap1[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [3];
assign \w_pma_adapt_dfe_fltap1[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [4];
assign \w_pma_adapt_dfe_fltap1[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus [5];

assign \w_pma_adapt_dfe_fltap2[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [0];
assign \w_pma_adapt_dfe_fltap2[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [1];
assign \w_pma_adapt_dfe_fltap2[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [2];
assign \w_pma_adapt_dfe_fltap2[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [3];
assign \w_pma_adapt_dfe_fltap2[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [4];
assign \w_pma_adapt_dfe_fltap2[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus [5];

assign \w_pma_adapt_dfe_fltap3[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [0];
assign \w_pma_adapt_dfe_fltap3[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [1];
assign \w_pma_adapt_dfe_fltap3[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [2];
assign \w_pma_adapt_dfe_fltap3[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [3];
assign \w_pma_adapt_dfe_fltap3[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [4];
assign \w_pma_adapt_dfe_fltap3[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus [5];

assign \w_pma_adapt_dfe_fltap4[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [0];
assign \w_pma_adapt_dfe_fltap4[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [1];
assign \w_pma_adapt_dfe_fltap4[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [2];
assign \w_pma_adapt_dfe_fltap4[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [3];
assign \w_pma_adapt_dfe_fltap4[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [4];
assign \w_pma_adapt_dfe_fltap4[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus [5];

assign \w_pma_adapt_dfe_fltap_position[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [0];
assign \w_pma_adapt_dfe_fltap_position[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [1];
assign \w_pma_adapt_dfe_fltap_position[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [2];
assign \w_pma_adapt_dfe_fltap_position[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [3];
assign \w_pma_adapt_dfe_fltap_position[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [4];
assign \w_pma_adapt_dfe_fltap_position[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus [5];

assign \w_pma_adapt_dfe_fxtap1[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [0];
assign \w_pma_adapt_dfe_fxtap1[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [1];
assign \w_pma_adapt_dfe_fxtap1[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [2];
assign \w_pma_adapt_dfe_fxtap1[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [3];
assign \w_pma_adapt_dfe_fxtap1[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [4];
assign \w_pma_adapt_dfe_fxtap1[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [5];
assign \w_pma_adapt_dfe_fxtap1[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus [6];

assign \w_pma_adapt_dfe_fxtap2[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [0];
assign \w_pma_adapt_dfe_fxtap2[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [1];
assign \w_pma_adapt_dfe_fxtap2[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [2];
assign \w_pma_adapt_dfe_fxtap2[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [3];
assign \w_pma_adapt_dfe_fxtap2[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [4];
assign \w_pma_adapt_dfe_fxtap2[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [5];
assign \w_pma_adapt_dfe_fxtap2[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus [6];

assign \w_pma_adapt_dfe_fxtap3[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [0];
assign \w_pma_adapt_dfe_fxtap3[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [1];
assign \w_pma_adapt_dfe_fxtap3[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [2];
assign \w_pma_adapt_dfe_fxtap3[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [3];
assign \w_pma_adapt_dfe_fxtap3[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [4];
assign \w_pma_adapt_dfe_fxtap3[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [5];
assign \w_pma_adapt_dfe_fxtap3[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus [6];

assign \w_pma_adapt_dfe_fxtap4[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [0];
assign \w_pma_adapt_dfe_fxtap4[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [1];
assign \w_pma_adapt_dfe_fxtap4[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [2];
assign \w_pma_adapt_dfe_fxtap4[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [3];
assign \w_pma_adapt_dfe_fxtap4[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [4];
assign \w_pma_adapt_dfe_fxtap4[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus [5];

assign \w_pma_adapt_dfe_fxtap5[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [0];
assign \w_pma_adapt_dfe_fxtap5[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [1];
assign \w_pma_adapt_dfe_fxtap5[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [2];
assign \w_pma_adapt_dfe_fxtap5[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [3];
assign \w_pma_adapt_dfe_fxtap5[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [4];
assign \w_pma_adapt_dfe_fxtap5[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus [5];

assign \w_pma_adapt_dfe_fxtap6[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus [0];
assign \w_pma_adapt_dfe_fxtap6[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus [1];
assign \w_pma_adapt_dfe_fxtap6[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus [2];
assign \w_pma_adapt_dfe_fxtap6[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus [3];
assign \w_pma_adapt_dfe_fxtap6[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus [4];

assign \w_pma_adapt_dfe_fxtap7[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus [0];
assign \w_pma_adapt_dfe_fxtap7[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus [1];
assign \w_pma_adapt_dfe_fxtap7[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus [2];
assign \w_pma_adapt_dfe_fxtap7[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus [3];
assign \w_pma_adapt_dfe_fxtap7[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus [4];

assign \w_pma_adapt_odi_vref[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus [0];
assign \w_pma_adapt_odi_vref[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus [1];
assign \w_pma_adapt_odi_vref[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus [2];
assign \w_pma_adapt_odi_vref[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus [3];
assign \w_pma_adapt_odi_vref[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus [4];

assign \w_pma_adapt_vga_sel[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [0];
assign \w_pma_adapt_vga_sel[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [1];
assign \w_pma_adapt_vga_sel[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [2];
assign \w_pma_adapt_vga_sel[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [3];
assign \w_pma_adapt_vga_sel[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [4];
assign \w_pma_adapt_vga_sel[5]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [5];
assign \w_pma_adapt_vga_sel[6]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus [6];

assign \w_pma_adapt_vref_sel[0]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus [0];
assign \w_pma_adapt_vref_sel[1]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus [1];
assign \w_pma_adapt_vref_sel[2]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus [2];
assign \w_pma_adapt_vref_sel[3]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus [3];
assign \w_pma_adapt_vref_sel[4]  = \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus [4];

twentynm_hssi_pma_tx_buf \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.bsmode(gnd),
	.bsoeb(gnd),
	.bstxn_in(gnd),
	.bstxp_in(gnd),
	.clk0_tx(w_pma_cgb_hifreqclkp),
	.clk180_tx(w_pma_cgb_hifreqclkn),
	.clk_dcd(\w_pma_cgb_cpulse_out_bus[0] ),
	.clksn(w_pma_tx_ser_ckdrvp),
	.clksp(w_pma_tx_ser_ckdrvn),
	.cr_rdynamic_sw(),
	.oe(w_pma_tx_ser_oe),
	.oeb(w_pma_tx_ser_oeb),
	.oo(w_pma_tx_ser_oo),
	.oob(w_pma_tx_ser_oob),
	.pcie_sw_master(\w_pma_cgb_pcie_sw_master[1] ),
	.rx_det_clk(w_pma_cdr_refclk_rx_det_clk),
	.rx_n_bidir_in(gnd),
	.rx_p_bidir_in(in_rx_p),
	.s_lpbk_b(in_rs_lpbk_b),
	.tx_det_rx(in_tx_det_rx),
	.tx_elec_idle(in_tx_elec_idle),
	.tx_qpi_pulldn(in_tx_qpi_pulldn),
	.tx_qpi_pullup(in_tx_qpi_pullup),
	.tx_rlpbk(w_cdr_pll_tx_rlpbk),
	.vrlpbkn(w_cdr_pll_rlpbkn),
	.vrlpbkn_1t(w_cdr_pll_rlpbkdn),
	.vrlpbkp(w_cdr_pll_rlpbkp),
	.vrlpbkp_1t(w_cdr_pll_rlpbkdp),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.i_coeff({in_i_coeff[17],in_i_coeff[16],in_i_coeff[15],in_i_coeff[14],in_i_coeff[13],in_i_coeff[12],in_i_coeff[11],in_i_coeff[10],in_i_coeff[9],in_i_coeff[8],in_i_coeff[7],in_i_coeff[6],in_i_coeff[5],in_i_coeff[4],in_i_coeff[3],in_i_coeff[2],in_i_coeff[1],in_i_coeff[0]}),
	.tx50({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.blockselect(out_blockselect_pma_tx_buf),
	.ckn(w_pma_tx_buf_ckn),
	.ckp(w_pma_tx_buf_ckp),
	.dcd_out1(),
	.dcd_out2(),
	.dcd_out_ready(),
	.lbvon(w_pma_tx_buf_lbvon),
	.lbvop(w_pma_tx_buf_lbvop),
	.rx_detect_valid(out_rx_detect_valid),
	.rx_found(out_rx_found),
	.rx_found_pcie_spl_test(),
	.sel_vreg(),
	.spl_clk_test(),
	.vlptxn(),
	.vlptxp(),
	.von(),
	.vop(out_tx_p),
	.atbsel(\gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_ATBSEL_bus ),
	.avmmreaddata(\gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf_AVMMREADDATA_bus ),
	.detect_on(),
	.tx_dftout());
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .calibration_en = "false";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .calibration_resistor_value = "res_setting0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .cdr_cp_calibration_en = "cdr_cp_cal_disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .chgpmp_current_dn_trim = "cp_current_trimming_dn_setting0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .chgpmp_current_up_trim = "cp_current_trimming_up_setting0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .chgpmp_dn_trim_double = "normal_dn_trim_current";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .chgpmp_up_trim_double = "normal_up_trim_current";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .compensation_driver_en = "disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .compensation_en = "enable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .cpen_ctrl = "cp_l0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .dcd_clk_div_ctrl = "dcd_ck_div128";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .dcd_detection_en = "enable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .dft_sel = "dft_disabled";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_bandwidth = "dcc_bw_12";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_bandwidth_dn = "dcd_bw_dn_0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_mode_ctrl = "dcc_disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_reference1 = "dcc_ref1_3";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_reference2 = "dcc_ref2_3";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_correction_reset_n = "reset_n";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_cp_comp_en = "cp_comp_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_detector_cp_cal = "dcd_cp_cal_disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_detector_sa_cal = "dcd_sa_cal_disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_input_polarity = "dcc_input_pos";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_setting = "dcc_t32";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .duty_cycle_setting_aux = "dcc2_t32";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .enable_idle_tx_channel_support = "false";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .jtag_drv_sel = "drv1";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .jtag_lp = "lp_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .link = "sr";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .link_tx = "sr";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .low_power_en = "disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .lst = "atb_disabled";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .mcgb_location_for_pcie = 4'b0000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .optimal = "false";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pm_speed_grade = "e2";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .power_rail_eht = 0;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .power_rail_et = 0;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_sign_1st_post_tap = "fir_post_1t_neg";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_sign_2nd_post_tap = "fir_post_2t_neg";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_sign_pre_tap_1t = "fir_pre_1t_neg";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_sign_pre_tap_2t = "fir_pre_2t_neg";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_switching_ctrl_1st_post_tap = 6'b000000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_switching_ctrl_2nd_post_tap = 4'b0000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_switching_ctrl_pre_tap_1t = 5'b00000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .pre_emp_switching_ctrl_pre_tap_2t = 3'b000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .prot_mode = "basic_tx";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .res_cal_local = "non_local";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .rx_det = "mode_0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .rx_det_output_sel = "rx_det_pcie_out";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .rx_det_pdb = "rx_det_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .sense_amp_offset_cal_curr_n = "sa_os_cal_in_0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .sense_amp_offset_cal_curr_p = 5'b00000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .ser_powerdown = "normal_ser_on";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .slew_rate_ctrl = "slew_r7";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .swing_level = "lv";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .term_code = "rterm_code7";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .term_n_tune = "rterm_n0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .term_p_tune = "rterm_p0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .term_sel = "r_r1";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .tri_driver = "tri_driver_disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .tx_powerdown = "normal_tx_on";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_dcd_cal = "uc_dcd_cal_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_dcd_cal_status = "uc_dcd_cal_notdone";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_gen3 = "gen3_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_gen4 = "gen4_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_skew_cal = "uc_skew_cal_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_skew_cal_status = "uc_skew_cal_notdone";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_txvod_cal = "uc_tx_vod_cal_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_txvod_cal_cont = "uc_tx_vod_cal_cont_off";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_txvod_cal_status = "uc_tx_vod_cal_notdone";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .uc_vcc_setting = "vcc_setting0";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .user_fir_coeff_ctrl_sel = "ram_ctl";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .vod_output_swing_ctrl = 5'b00000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .vreg_output = "vccdreg_nominal";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_analog_mode = "user_custom";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_bonding_mode = "x1_non_bonded";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_calibration_en = "false";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_clock_divider_ratio = 4'b0100;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_datawidth = 8'b00001010;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_gt_enabled = "disable";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_initial_settings = "true";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_optimal = "false";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_pma_tx_divclk_hz = 32'b00000111011100110101100101000000;
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_prot_mode = "basic_tx";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_swing_level = "lv";
defparam \gen_twentynm_hssi_pma_tx_buf.inst_twentynm_hssi_pma_tx_buf .xtx_path_tx_pll_clk_hz = "156250000";

twentynm_hssi_pma_tx_ser \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.bitslipstate(w_pma_cgb_bitslipstate),
	.cpulse(\w_pma_cgb_cpulse_out_bus[1] ),
	.hfclkn(\w_pma_cgb_cpulse_out_bus[4] ),
	.hfclkp(\w_pma_cgb_cpulse_out_bus[5] ),
	.lfclk(\w_pma_cgb_cpulse_out_bus[3] ),
	.lfclk2(\w_pma_cgb_cpulse_out_bus[2] ),
	.paraclk(\w_pma_cgb_cpulse_out_bus[0] ),
	.rser_div2(w_pma_cgb_div2),
	.rser_div4(w_pma_cgb_div4),
	.rser_div5(w_pma_cgb_div5),
	.rst_n(w_pma_cgb_rstb),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.data({in_tx_data[63],in_tx_data[62],in_tx_data[61],in_tx_data[60],in_tx_data[59],in_tx_data[58],in_tx_data[57],in_tx_data[56],in_tx_data[55],in_tx_data[54],in_tx_data[53],in_tx_data[52],in_tx_data[51],in_tx_data[50],in_tx_data[49],in_tx_data[48],in_tx_data[47],in_tx_data[46],in_tx_data[45],in_tx_data[44],in_tx_data[43],in_tx_data[42],in_tx_data[41],in_tx_data[40],in_tx_data[39],
in_tx_data[38],in_tx_data[37],in_tx_data[36],in_tx_data[35],in_tx_data[34],in_tx_data[33],in_tx_data[32],in_tx_data[31],in_tx_data[30],in_tx_data[29],in_tx_data[28],in_tx_data[27],in_tx_data[26],in_tx_data[25],in_tx_data[24],in_tx_data[23],in_tx_data[22],in_tx_data[21],in_tx_data[20],in_tx_data[19],in_tx_data[18],in_tx_data[17],in_tx_data[16],in_tx_data[15],in_tx_data[14],
in_tx_data[13],in_tx_data[12],in_tx_data[11],in_tx_data[10],in_tx_data[9],in_tx_data[8],in_tx_data[7],in_tx_data[6],in_tx_data[5],in_tx_data[4],in_tx_data[3],in_tx_data[2],in_tx_data[1],in_tx_data[0]}),
	.blockselect(out_blockselect_pma_tx_ser),
	.ckdrvn(w_pma_tx_ser_ckdrvn),
	.ckdrvp(w_pma_tx_ser_ckdrvp),
	.clk_divtx(out_iqtxrxclk_out1),
	.clk_divtx_user(out_clkdiv_tx_user),
	.oe(w_pma_tx_ser_oe),
	.oeb(w_pma_tx_ser_oeb),
	.oo(w_pma_tx_ser_oo),
	.oob(w_pma_tx_ser_oob),
	.avmmreaddata(\gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser_AVMMREADDATA_bus ));
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .bonding_mode = "x1_non_bonded";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .clk_divtx_deskew = "deskew_delay8";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .control_clk_divtx = "no_dft_control_clkdivtx";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .duty_cycle_correction_mode_ctrl = "dcc_disable";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .prot_mode = "basic_tx";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .ser_clk_divtx_user_sel = "divtx_user_off";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .ser_clk_mon = "disable_clk_mon";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .ser_powerdown = "normal_poweron_ser";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_tx_ser.inst_twentynm_hssi_pma_tx_ser .sup_mode = "user_mode";

twentynm_hssi_pma_tx_cgb \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.ckdccn(w_pma_tx_buf_ckn),
	.ckdccp(w_pma_tx_buf_ckp),
	.clk_cdr_b(gnd),
	.clk_cdr_direct(w_cdr_pll_clk0_pfd),
	.clk_cdr_t(gnd),
	.clk_fpll_b(in_clk_fpll_b),
	.clk_fpll_t(gnd),
	.clk_lc_b(gnd),
	.clk_lc_hs(gnd),
	.clk_lc_t(gnd),
	.clkb_cdr_b(gnd),
	.clkb_cdr_direct(w_cdr_pll_clk180_pfd),
	.clkb_cdr_t(gnd),
	.clkb_fpll_b(gnd),
	.clkb_fpll_t(gnd),
	.clkb_lc_b(gnd),
	.clkb_lc_hs(gnd),
	.clkb_lc_t(gnd),
	.tx_bitslip(in_tx_bitslip),
	.tx_bonding_rstb(in_tx_bonding_rstb),
	.tx_pma_rstb(in_tx_pma_rstb),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.cpulse_x6_dn_bus({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cpulse_x6_up_bus({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cpulse_xn_dn_bus({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cpulse_xn_up_bus({gnd,gnd,gnd,gnd,gnd,gnd}),
	.pcie_sw({in_pcie_sw[1],in_pcie_sw[0]}),
	.pcie_sw_done_master({gnd,gnd}),
	.bitslipstate(w_pma_cgb_bitslipstate),
	.blockselect(out_blockselect_pma_cgb),
	.div2(w_pma_cgb_div2),
	.div4(w_pma_cgb_div4),
	.div5(w_pma_cgb_div5),
	.hifreqclkn(w_pma_cgb_hifreqclkn),
	.hifreqclkp(w_pma_cgb_hifreqclkp),
	.rstb(w_pma_cgb_rstb),
	.avmmreaddata(\gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_AVMMREADDATA_bus ),
	.cpulse_out_bus(\gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_CPULSE_OUT_BUS_bus ),
	.pcie_sw_done(\gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_DONE_bus ),
	.pcie_sw_master(\gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb_PCIE_SW_MASTER_bus ));
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .bitslip_enable = "disable_bitslip";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .bonding_mode = "x1_non_bonded";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .bonding_reset_enable = "disallow_bonding_reset";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .cgb_power_down = "normal_cgb";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .dprio_cgb_vreg_boost = "no_voltage_boost";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .input_select_gen3 = "unused";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .input_select_x1 = "fpll_bot";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .input_select_xn = "unused";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .observe_cgb_clocks = "observe_nothing";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .pcie_gen3_bitwidth = "pciegen3_wide";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .prot_mode = "basic_tx";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .scratch0_x1_clock_src = "fpll_bot";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .scratch1_x1_clock_src = "unused";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .scratch2_x1_clock_src = "unused";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .scratch3_x1_clock_src = "unused";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .select_done_master_or_slave = "choose_slave_pcie_sw_done";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .ser_mode = "ten_bit";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .ser_powerdown = "normal_poweron_ser";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .tx_ucontrol_en = "disable";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .tx_ucontrol_pcie = "gen1";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .tx_ucontrol_reset = "disable";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .vccdreg_output = "vccdreg_nominal";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .x1_clock_source_sel = "cdr_txpll_t";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .x1_div_m_sel = "divby4";
defparam \gen_twentynm_hssi_pma_tx_cgb.inst_twentynm_hssi_pma_tx_cgb .xn_clock_source_sel = "sel_xn_up";

twentynm_hssi_pma_rx_deser \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser (
	.adapt_en(\w_pma_adapt_odi_vref[0] ),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.bitslip(in_rx_bitslip),
	.clk0(w_cdr_pll_clk0_des),
	.clk0_odi(w_pma_rx_odi_clk0_eye),
	.clk180(w_cdr_pll_clk180_des),
	.clk180_odi(w_pma_rx_odi_clk180_eye),
	.clk270(),
	.clk90(),
	.clklow(out_clklow),
	.deven(w_cdr_pll_deven_des),
	.deven_odi(w_pma_rx_odi_de_eye),
	.devenb(w_cdr_pll_devenb_des),
	.devenb_odi(w_pma_rx_odi_deb_eye),
	.dodd(w_cdr_pll_dodd_des),
	.dodd_odi(w_pma_rx_odi_do_eye),
	.doddb(w_cdr_pll_doddb_des),
	.doddb_odi(w_pma_rx_odi_dob_eye),
	.error_even(w_cdr_pll_error_even_des),
	.error_evenb(w_cdr_pll_error_evenb_des),
	.error_odd(w_cdr_pll_error_odd_des),
	.error_oddb(w_cdr_pll_error_oddb_des),
	.fref(out_fref),
	.odi_en(w_pma_rx_odi_odi_en),
	.pfdmode_lock(out_pfdmode_lock),
	.rst_n(in_rx_pma_rstb),
	.tdr_en(),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.pcie_sw({in_pcie_sw[1],in_pcie_sw[0]}),
	.adapt_clk(w_pma_rx_deser_adapt_clk),
	.blockselect(out_blockselect_pma_rx_deser),
	.clkdiv(out_clkdiv_rx),
	.clkdiv_user(out_clkdiv_rx_user),
	.clkdivrx_rx(w_pma_rx_deser_clkdivrx_rx),
	.odi_clkout(),
	.avmmreaddata(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_AVMMREADDATA_bus ),
	.data(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DATA_bus ),
	.dout(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_DOUT_bus ),
	.error_deser(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ERROR_DESER_bus ),
	.odi_dout(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_ODI_DOUT_bus ),
	.pcie_sw_ret(\gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser_PCIE_SW_RET_bus ),
	.tstmx_deser());
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .bitslip_bypass = "bs_bypass_no";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .clkdiv_source = "vco_bypass_normal";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .clkdivrx_user_mode = "clkdivrx_user_disabled";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .deser_factor = 10;
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .deser_powerdown = "deser_power_up";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .force_adaptation_outputs = "normal_outputs";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .force_clkdiv_for_testing = "normal_clkdiv";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .pcie_gen = "non_pcie";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .pcie_gen_bitwidth = "pcie_gen3_32b";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .rst_n_adapt_odi = "no_rst_adapt_odi";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .sdclk_enable = "false";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_rx_deser.inst_twentynm_hssi_pma_rx_deser .tdr_mode = "select_bbpd_data";

twentynm_hssi_pma_rx_buf \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk_divrx(w_pma_rx_deser_clkdivrx_rx),
	.lpbkn(w_pma_tx_buf_lbvon),
	.lpbkp(w_pma_tx_buf_lbvop),
	.rx_qpi_pulldn(in_rx_qpi_pulldn),
	.rx_rstn(in_rx_pma_rstb),
	.rxn(gnd),
	.rxp(in_rx_p),
	.s_lpbk_b(in_rs_lpbk_b),
	.vga_cm_bidir_in(),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.rx_sel_b50({gnd,gnd,gnd,gnd,gnd,gnd}),
	.vcz({\w_pma_adapt_ctle_acgain_4s[27] ,\w_pma_adapt_ctle_acgain_4s[26] ,\w_pma_adapt_ctle_acgain_4s[25] ,\w_pma_adapt_ctle_acgain_4s[24] ,\w_pma_adapt_ctle_acgain_4s[23] ,\w_pma_adapt_ctle_acgain_4s[22] ,\w_pma_adapt_ctle_acgain_4s[21] ,\w_pma_adapt_ctle_acgain_4s[20] ,
\w_pma_adapt_ctle_acgain_4s[19] ,\w_pma_adapt_ctle_acgain_4s[18] ,\w_pma_adapt_ctle_acgain_4s[17] ,\w_pma_adapt_ctle_acgain_4s[16] ,\w_pma_adapt_ctle_acgain_4s[15] ,\w_pma_adapt_ctle_acgain_4s[14] ,\w_pma_adapt_ctle_acgain_4s[13] ,\w_pma_adapt_ctle_acgain_4s[12] ,
\w_pma_adapt_ctle_acgain_4s[11] ,\w_pma_adapt_ctle_acgain_4s[10] ,\w_pma_adapt_ctle_acgain_4s[9] ,\w_pma_adapt_ctle_acgain_4s[8] ,\w_pma_adapt_ctle_acgain_4s[7] ,\w_pma_adapt_ctle_acgain_4s[6] ,\w_pma_adapt_ctle_acgain_4s[5] ,\w_pma_adapt_ctle_acgain_4s[4] ,
\w_pma_adapt_ctle_acgain_4s[3] ,\w_pma_adapt_ctle_acgain_4s[2] ,\w_pma_adapt_ctle_acgain_4s[1] ,\w_pma_adapt_ctle_acgain_4s[0] }),
	.vds_eqz_s1_set({\w_pma_adapt_ctle_eqz_1s_sel[14] ,\w_pma_adapt_ctle_eqz_1s_sel[13] ,\w_pma_adapt_ctle_eqz_1s_sel[12] ,\w_pma_adapt_ctle_eqz_1s_sel[11] ,\w_pma_adapt_ctle_eqz_1s_sel[10] ,\w_pma_adapt_ctle_eqz_1s_sel[9] ,\w_pma_adapt_ctle_eqz_1s_sel[8] ,
\w_pma_adapt_ctle_eqz_1s_sel[7] ,\w_pma_adapt_ctle_eqz_1s_sel[6] ,\w_pma_adapt_ctle_eqz_1s_sel[5] ,\w_pma_adapt_ctle_eqz_1s_sel[4] ,\w_pma_adapt_ctle_eqz_1s_sel[3] ,\w_pma_adapt_ctle_eqz_1s_sel[2] ,\w_pma_adapt_ctle_eqz_1s_sel[1] ,\w_pma_adapt_ctle_eqz_1s_sel[0] }),
	.vds_lfeqz_czero({gnd,gnd}),
	.vds_lfeqz_fb_set({\w_pma_adapt_ctle_lfeq_fb_sel[6] ,\w_pma_adapt_ctle_lfeq_fb_sel[5] ,\w_pma_adapt_ctle_lfeq_fb_sel[4] ,\w_pma_adapt_ctle_lfeq_fb_sel[3] ,\w_pma_adapt_ctle_lfeq_fb_sel[2] ,\w_pma_adapt_ctle_lfeq_fb_sel[1] ,\w_pma_adapt_ctle_lfeq_fb_sel[0] }),
	.vds_vga_set({\w_pma_adapt_vga_sel[6] ,\w_pma_adapt_vga_sel[5] ,\w_pma_adapt_vga_sel[4] ,\w_pma_adapt_vga_sel[3] ,\w_pma_adapt_vga_sel[2] ,\w_pma_adapt_vga_sel[1] ,\w_pma_adapt_vga_sel[0] }),
	.blockselect(out_blockselect_pma_rx_buf),
	.inn(w_pma_rx_buf_inn),
	.inp(w_pma_rx_buf_inp),
	.outn(w_pma_rx_buf_outn),
	.outp(w_pma_rx_buf_outp),
	.pull_dn(w_pma_rx_buf_pull_dn),
	.rdlpbkn(w_pma_rx_buf_rdlpbkn),
	.rdlpbkp(w_pma_rx_buf_rdlpbkp),
	.rx_refclk(),
	.vga_cm_bidir_out(),
	.avmmreaddata(\gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf_AVMMREADDATA_bus ));
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .act_isource_disable = "isrc_en";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .bodybias_enable = "bodybias_en";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .bodybias_select = "bodybias_sel1";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .bypass_eqz_stages_234 = "bypass_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .cdrclk_to_cgb = "cdrclk_2cgb_dis";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .cgm_bias_disable = "cgmbias_en";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .diag_lp_en = "dlp_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .eq_bw_sel = "eq_bw_1";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .eq_dc_gain_trim = "no_dc_gain";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .input_vcm_sel = "high_vcm";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .iostandard = "hssi_diffio";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .lfeq_enable = "non_lfeq_mode";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .lfeq_zero_control = "lfeq_setting_2";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .link = "sr";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .link_rx = "sr";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .loopback_modes = "lpbk_disable";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .offset_cal_pd = "eqz1_en";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .offset_cancellation_coarse = "coarse_setting_00";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .offset_cancellation_ctrl = "volt_0mv";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .offset_cancellation_fine = "fine_setting_00";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .offset_pd = "oc_en";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .one_stage_enable = "non_s1_mode";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pdb_rx = "normal_rx_on";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pm_speed_grade = "e2";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pm_tx_rx_cvp_mode = "cvp_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pm_tx_rx_pcie_gen = "non_pcie";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pm_tx_rx_pcie_gen_bitwidth = "pcie_gen3_32b";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .pm_tx_rx_testmux_select = "setting0";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .power_mode_rx = "low_power";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .power_rail_eht = 0;
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .power_rail_er = 0;
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .qpi_enable = "non_qpi_mode";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .refclk_en = "disable";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .rx_atb_select = "atb_disable";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .rx_refclk_divider = "bypass_divider";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .rx_sel_bias_source = "bias_vcmdrv";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .rx_vga_oc_en = "vga_cal_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .term_sel = "r_r1";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .term_tri_enable = "disable_tri";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .vccela_supply_voltage = "vccela_1p1v";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .vcm_current_add = "vcm_current_default";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .vcm_sel = "vcm_setting_10";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .vga_bandwidth_select = "vga_bw_1";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_analog_mode = "user_custom";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_datawidth = 8'b00001010;
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_gt_enabled = "disable";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_initial_settings = "true";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_jtag_hys = "hys_increase_disable";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_jtag_lp = "lp_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_pma_rx_divclk_hz = 32'b00000111011100110101100101000000;
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_uc_cal_enable = "rx_cal_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_uc_cru_rstb = "cdr_lf_reset_off";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_uc_pcie_sw = "uc_pcie_gen1";
defparam \gen_twentynm_hssi_pma_rx_buf.inst_twentynm_hssi_pma_rx_buf .xrx_path_uc_rx_rstb = "rx_reset_on";

twentynm_hssi_pma_rx_sd \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk(w_pma_rx_deser_clkdivrx_rx),
	.qpi(w_pma_rx_buf_pull_dn),
	.rstn_sd(in_rx_pma_rstb),
	.s_lpbk_b(in_rs_lpbk_b),
	.vin(w_pma_rx_buf_inn),
	.vip(w_pma_rx_buf_inp),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.blockselect(out_blockselect_pma_rx_sd),
	.sd(out_sd),
	.avmmreaddata(\gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd_AVMMREADDATA_bus ));
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .link = "sr";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .sd_output_off = 1;
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .sd_output_on = 15;
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .sd_pdb = "sd_off";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .sd_threshold = "sdlv_3";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_rx_sd.inst_twentynm_hssi_pma_rx_sd .sup_mode = "user_mode";

twentynm_hssi_pma_rx_odi \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk0(w_cdr_pll_clk0_odi),
	.clk180(w_cdr_pll_clk180_odi),
	.clk270(w_cdr_pll_clk270_odi),
	.clk90(w_cdr_pll_clk90_odi),
	.it50u(),
	.it50u2(),
	.it50u4(),
	.odi_dft_clr(in_eye_monitor[3]),
	.odi_latch_clk(in_eye_monitor[1]),
	.odi_shift_clk(in_eye_monitor[0]),
	.odi_shift_in(in_eye_monitor[2]),
	.rx_n(w_pma_rx_buf_inn),
	.rx_p(w_pma_rx_buf_inp),
	.rxn_sum(w_pma_rx_buf_outn),
	.rxp_sum(w_pma_rx_buf_outp),
	.spec_vrefh(w_pma_rx_dfe_spec_vrefh),
	.spec_vrefl(w_pma_rx_dfe_spec_vrefl),
	.vcm_vref(gnd),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.odi_atb_sel(),
	.vertical_fb({\w_pma_adapt_odi_vref[4] ,\w_pma_adapt_odi_vref[3] ,\w_pma_adapt_odi_vref[2] ,\w_pma_adapt_odi_vref[1] ,gnd}),
	.atb0(\gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi~atb0 ),
	.atb1(),
	.blockselect(out_blockselect_pma_rx_odi),
	.clk0_eye(w_pma_rx_odi_clk0_eye),
	.clk0_eye_lb(w_pma_rx_odi_clk0_eye_lb),
	.clk180_eye(w_pma_rx_odi_clk180_eye),
	.clk180_eye_lb(w_pma_rx_odi_clk180_eye_lb),
	.de_eye(w_pma_rx_odi_de_eye),
	.deb_eye(w_pma_rx_odi_deb_eye),
	.do_eye(w_pma_rx_odi_do_eye),
	.dob_eye(w_pma_rx_odi_dob_eye),
	.odi_en(w_pma_rx_odi_odi_en),
	.tdr_en(),
	.vref_sel_out(),
	.avmmreaddata(\gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi_AVMMREADDATA_bus ),
	.odi_oc_tstmx());
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .clk_dcd_bypass = "no_bypass";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .enable_odi = "power_down_eye";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .invert_dfe_vref = "no_inversion";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .monitor_bw_sel = "bw_1";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .oc_sa_c0 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .oc_sa_c180 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .phase_steps_64_vs_128 = "phase_steps_64";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .phase_steps_sel = "step40";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .sel_oc_en = "off_canc_disable";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .step_ctrl_sel = "dprio_mode";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .v_vert_sel = "plus";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .v_vert_threshold_scaling = "scale_3";
defparam \gen_twentynm_hssi_pma_rx_odi.inst_twentynm_hssi_pma_rx_odi .vert_threshold = "vert_0";

twentynm_hssi_pma_rx_dfe \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe (
	.adapt_en(w_pma_adapt_dfe_adapt_en),
	.adp_clk(w_pma_adapt_dfe_adp_clk),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk0(w_cdr_pll_clk0_pd),
	.clk180(w_cdr_pll_clk180_pd),
	.clk270(w_cdr_pll_clk270_pd),
	.clk90(w_cdr_pll_clk90_pd),
	.dfe_fltap1_sgn(w_pma_adapt_dfe_fltap1_sgn),
	.dfe_fltap2_sgn(w_pma_adapt_dfe_fltap2_sgn),
	.dfe_fltap3_sgn(w_pma_adapt_dfe_fltap3_sgn),
	.dfe_fltap4_sgn(w_pma_adapt_dfe_fltap4_sgn),
	.dfe_fltap_bypdeser(w_pma_adapt_dfe_fltap_bypdeser),
	.dfe_fxtap2_sgn(w_pma_adapt_dfe_fxtap2_sgn),
	.dfe_fxtap3_sgn(w_pma_adapt_dfe_fxtap3_sgn),
	.dfe_fxtap4_sgn(w_pma_adapt_dfe_fxtap4_sgn),
	.dfe_fxtap5_sgn(w_pma_adapt_dfe_fxtap5_sgn),
	.dfe_fxtap6_sgn(w_pma_adapt_dfe_fxtap6_sgn),
	.dfe_fxtap7_sgn(w_pma_adapt_dfe_fxtap7_sgn),
	.dfe_rstn(in_rx_pma_rstb),
	.dfe_spec_disable(w_pma_adapt_dfe_spec_disable),
	.dfe_spec_sgn_sel(w_pma_adapt_dfe_spec_sign_sel),
	.dfe_vref_sgn_sel(w_pma_adapt_dfe_vref_sign_sel),
	.rxn(w_pma_rx_buf_outn),
	.rxp(w_pma_rx_buf_outp),
	.vga_vcm(gnd),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.dfe_fltap1_coeff({\w_pma_adapt_dfe_fltap1[5] ,\w_pma_adapt_dfe_fltap1[4] ,\w_pma_adapt_dfe_fltap1[3] ,\w_pma_adapt_dfe_fltap1[2] ,\w_pma_adapt_dfe_fltap1[1] ,\w_pma_adapt_dfe_fltap1[0] }),
	.dfe_fltap2_coeff({\w_pma_adapt_dfe_fltap2[5] ,\w_pma_adapt_dfe_fltap2[4] ,\w_pma_adapt_dfe_fltap2[3] ,\w_pma_adapt_dfe_fltap2[2] ,\w_pma_adapt_dfe_fltap2[1] ,\w_pma_adapt_dfe_fltap2[0] }),
	.dfe_fltap3_coeff({\w_pma_adapt_dfe_fltap3[5] ,\w_pma_adapt_dfe_fltap3[4] ,\w_pma_adapt_dfe_fltap3[3] ,\w_pma_adapt_dfe_fltap3[2] ,\w_pma_adapt_dfe_fltap3[1] ,\w_pma_adapt_dfe_fltap3[0] }),
	.dfe_fltap4_coeff({\w_pma_adapt_dfe_fltap4[5] ,\w_pma_adapt_dfe_fltap4[4] ,\w_pma_adapt_dfe_fltap4[3] ,\w_pma_adapt_dfe_fltap4[2] ,\w_pma_adapt_dfe_fltap4[1] ,\w_pma_adapt_dfe_fltap4[0] }),
	.dfe_fltap_position({\w_pma_adapt_dfe_fltap_position[5] ,\w_pma_adapt_dfe_fltap_position[4] ,\w_pma_adapt_dfe_fltap_position[3] ,\w_pma_adapt_dfe_fltap_position[2] ,\w_pma_adapt_dfe_fltap_position[1] ,\w_pma_adapt_dfe_fltap_position[0] }),
	.dfe_fxtap1_coeff({\w_pma_adapt_dfe_fxtap1[6] ,\w_pma_adapt_dfe_fxtap1[5] ,\w_pma_adapt_dfe_fxtap1[4] ,\w_pma_adapt_dfe_fxtap1[3] ,\w_pma_adapt_dfe_fxtap1[2] ,\w_pma_adapt_dfe_fxtap1[1] ,\w_pma_adapt_dfe_fxtap1[0] }),
	.dfe_fxtap2_coeff({\w_pma_adapt_dfe_fxtap2[6] ,\w_pma_adapt_dfe_fxtap2[5] ,\w_pma_adapt_dfe_fxtap2[4] ,\w_pma_adapt_dfe_fxtap2[3] ,\w_pma_adapt_dfe_fxtap2[2] ,\w_pma_adapt_dfe_fxtap2[1] ,\w_pma_adapt_dfe_fxtap2[0] }),
	.dfe_fxtap3_coeff({\w_pma_adapt_dfe_fxtap3[6] ,\w_pma_adapt_dfe_fxtap3[5] ,\w_pma_adapt_dfe_fxtap3[4] ,\w_pma_adapt_dfe_fxtap3[3] ,\w_pma_adapt_dfe_fxtap3[2] ,\w_pma_adapt_dfe_fxtap3[1] ,\w_pma_adapt_dfe_fxtap3[0] }),
	.dfe_fxtap4_coeff({\w_pma_adapt_dfe_fxtap4[5] ,\w_pma_adapt_dfe_fxtap4[4] ,\w_pma_adapt_dfe_fxtap4[3] ,\w_pma_adapt_dfe_fxtap4[2] ,\w_pma_adapt_dfe_fxtap4[1] ,\w_pma_adapt_dfe_fxtap4[0] }),
	.dfe_fxtap5_coeff({\w_pma_adapt_dfe_fxtap5[5] ,\w_pma_adapt_dfe_fxtap5[4] ,\w_pma_adapt_dfe_fxtap5[3] ,\w_pma_adapt_dfe_fxtap5[2] ,\w_pma_adapt_dfe_fxtap5[1] ,\w_pma_adapt_dfe_fxtap5[0] }),
	.dfe_fxtap6_coeff({\w_pma_adapt_dfe_fxtap6[4] ,\w_pma_adapt_dfe_fxtap6[3] ,\w_pma_adapt_dfe_fxtap6[2] ,\w_pma_adapt_dfe_fxtap6[1] ,\w_pma_adapt_dfe_fxtap6[0] }),
	.dfe_fxtap7_coeff({\w_pma_adapt_dfe_fxtap7[4] ,\w_pma_adapt_dfe_fxtap7[3] ,\w_pma_adapt_dfe_fxtap7[2] ,\w_pma_adapt_dfe_fxtap7[1] ,\w_pma_adapt_dfe_fxtap7[0] }),
	.vref_level_coeff({\w_pma_adapt_vref_sel[4] ,\w_pma_adapt_vref_sel[3] ,\w_pma_adapt_vref_sel[2] ,\w_pma_adapt_vref_sel[1] ,\w_pma_adapt_vref_sel[0] }),
	.blockselect(out_blockselect_pma_rx_dfe),
	.clk0_bbpd(w_pma_rx_dfe_clk0_bbpd),
	.clk180_bbpd(w_pma_rx_dfe_clk180_bbpd),
	.clk270_bbpd(w_pma_rx_dfe_clk270_bbpd),
	.clk90_bbpd(w_pma_rx_dfe_clk90_bbpd),
	.deven(w_pma_rx_dfe_deven),
	.devenb(w_pma_rx_dfe_devenb),
	.dodd(w_pma_rx_dfe_dodd),
	.doddb(w_pma_rx_dfe_doddb),
	.edge270(w_pma_rx_dfe_edge270),
	.edge270b(w_pma_rx_dfe_edge270b),
	.edge90(w_pma_rx_dfe_edge90),
	.edge90b(w_pma_rx_dfe_edge90b),
	.err_ev(w_pma_rx_dfe_err_ev),
	.err_evb(w_pma_rx_dfe_err_evb),
	.err_od(w_pma_rx_dfe_err_od),
	.err_odb(w_pma_rx_dfe_err_odb),
	.spec_vrefh(w_pma_rx_dfe_spec_vrefh),
	.spec_vrefl(w_pma_rx_dfe_spec_vrefl),
	.avmmreaddata(\gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe_AVMMREADDATA_bus ),
	.dfe_oc_tstmx());
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .atb_select = "atb_disable";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .dft_en = "dft_disable";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_adp1 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_adp2 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_c270 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_c90 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_d0c0 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_d0c180 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_d1c0 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .oc_sa_d1c180 = 8'b00000000;
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .optimal = "false";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .pdb = "dfe_enable";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .pdb_fixedtap = "fixtap_dfe_powerdown";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .pdb_floattap = "floattap_dfe_powerdown";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .pdb_fxtap4t7 = "fxtap4t7_powerdown";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_fltapstep_dec = "fltap_step_no_dec";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_fltapstep_inc = "fltap_step_no_inc";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_fxtapstep_dec = "fxtap_step_no_dec";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_fxtapstep_inc = "fxtap_step_no_inc";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_oc_en = "off_canc_disable";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sel_probe_tstmx = "probe_tstmx_none";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .uc_rx_dfe_cal = "uc_rx_dfe_cal_off";
defparam \gen_twentynm_hssi_pma_rx_dfe.inst_twentynm_hssi_pma_rx_dfe .uc_rx_dfe_cal_status = "uc_rx_dfe_cal_notdone";

twentynm_hssi_pma_channel_pll \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll (
	.adapt_en(w_pma_adapt_dfe_adapt_en),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.clk0_bbpd(w_pma_rx_dfe_clk0_bbpd),
	.clk180_bbpd(w_pma_rx_dfe_clk180_bbpd),
	.clk270_bbpd(w_pma_rx_dfe_clk270_bbpd),
	.clk90_bbpd(w_pma_rx_dfe_clk90_bbpd),
	.deven(w_pma_rx_dfe_deven),
	.devenb(w_pma_rx_dfe_devenb),
	.dfe_test(gnd),
	.dodd(w_pma_rx_dfe_dodd),
	.doddb(w_pma_rx_dfe_doddb),
	.e270(w_pma_rx_dfe_edge270),
	.e270b(w_pma_rx_dfe_edge270b),
	.e90(w_pma_rx_dfe_edge90),
	.e90b(w_pma_rx_dfe_edge90b),
	.early_eios(in_early_eios),
	.error_even(w_pma_rx_dfe_err_ev),
	.error_evenb(w_pma_rx_dfe_err_evb),
	.error_odd(w_pma_rx_dfe_err_od),
	.error_oddb(w_pma_rx_dfe_err_odb),
	.fpll_test0(gnd),
	.fpll_test1(gnd),
	.ltd_b(in_ltd_b),
	.ltr(in_ltr),
	.odi_clk(w_pma_rx_odi_clk0_eye_lb),
	.odi_clkb(w_pma_rx_odi_clk180_eye_lb),
	.ppm_lock(in_ppm_lock),
	.refclk(w_pma_cdr_refclk_refclk),
	.rst_n(in_rx_pma_rstb),
	.rx_deser_pclk_test(w_pma_rx_deser_clkdivrx_rx),
	.rx_lpbkn(w_pma_rx_buf_rdlpbkn),
	.rx_lpbkp(w_pma_rx_buf_rdlpbkp),
	.rxp(in_rx_p),
	.sd(out_sd),
	.tx_ser_pclk_test(out_iqtxrxclk_out1),
	.atbsel(),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.iqtxrxclk({gnd,gnd,gnd,gnd,gnd,gnd}),
	.pcie_sw_ret({\w_pma_rx_deser_pcie_sw_ret[1] ,\w_pma_rx_deser_pcie_sw_ret[0] }),
	.blockselect(out_blockselect_cdr_pll),
	.cdr_cnt_done(),
	.cdr_lpbkdp(\gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll~O_CDR_LPBKDP ),
	.cdr_lpbkp(),
	.clk0_des(w_cdr_pll_clk0_des),
	.clk0_odi(w_cdr_pll_clk0_odi),
	.clk0_pd(w_cdr_pll_clk0_pd),
	.clk0_pfd(w_cdr_pll_clk0_pfd),
	.clk180_des(w_cdr_pll_clk180_des),
	.clk180_odi(w_cdr_pll_clk180_odi),
	.clk180_pd(w_cdr_pll_clk180_pd),
	.clk180_pfd(w_cdr_pll_clk180_pfd),
	.clk270_des(),
	.clk270_odi(w_cdr_pll_clk270_odi),
	.clk270_pd(w_cdr_pll_clk270_pd),
	.clk90_des(),
	.clk90_odi(w_cdr_pll_clk90_odi),
	.clk90_pd(w_cdr_pll_clk90_pd),
	.clklow(out_clklow),
	.deven_des(w_cdr_pll_deven_des),
	.devenb_des(w_cdr_pll_devenb_des),
	.dodd_des(w_cdr_pll_dodd_des),
	.doddb_des(w_cdr_pll_doddb_des),
	.error_even_des(w_cdr_pll_error_even_des),
	.error_evenb_des(w_cdr_pll_error_evenb_des),
	.error_odd_des(w_cdr_pll_error_odd_des),
	.error_oddb_des(w_cdr_pll_error_oddb_des),
	.fref(out_fref),
	.lock2ref(),
	.overrange(),
	.pfdmode_lock(out_pfdmode_lock),
	.rlpbkdn(w_cdr_pll_rlpbkdn),
	.rlpbkdp(w_cdr_pll_rlpbkdp),
	.rlpbkn(w_cdr_pll_rlpbkn),
	.rlpbkp(w_cdr_pll_rlpbkp),
	.rx_signal_ok(),
	.rxpll_lock(out_rxpll_lock),
	.tx_rlpbk(w_cdr_pll_tx_rlpbk),
	.underrange(),
	.von_lp(),
	.vop_lp(),
	.avmmreaddata(\gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll_AVMMREADDATA_bus ),
	.cdr_refclk_cal_out(),
	.cdr_vco_cal_out());
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .analog_mode = "user_custom";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .atb_select_control = "atb_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .auto_reset_on = "auto_reset_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .bandwidth_range_high = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .bandwidth_range_low = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .bbpd_data_pattern_filter_select = "bbpd_data_pat_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .bw_sel = "medium";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .cal_vco_count_length = "sel_8b_count";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .cdr_odi_select = "sel_cdr";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .cdr_phaselock_mode = "no_ignore_lock";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .cdr_powerdown_mode = "power_up";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .cgb_div = 1;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_dn_pd = "cp_current_pd_dn_setting4";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_dn_trim = "cp_current_trimming_dn_setting0";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_pd = "cp_current_pd_setting0";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_pfd = "cp_current_pfd_setting3";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_up_pd = "cp_current_pd_up_setting4";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_current_up_trim = "cp_current_trimming_up_setting0";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_dn_pd_trim_double = "normal_dn_trim_current";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_replicate = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_testmode = "cp_test_disable";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_up_pd_trim_double = "normal_up_trim_current";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .chgpmp_vccreg = "vreg_fw0";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .clklow_mux_select = "clklow_mux_cdr_fbclk";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .diag_loopback_enable = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .disable_up_dn = "true";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .enable_idle_rx_channel_support = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_max_cmu_out_freq = 36'b000000000000000000000000000000000001;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_max_m_counter = 36'b000000000000000000000000000000000001;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_max_pfd = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_max_ref = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_max_vco = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_min_gt_channel = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_min_pfd = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_min_ref = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .f_min_vco = "0 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .fb_select = "direct_fb";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .fref_clklow_div = 1;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .fref_mux_select = "fref_mux_cdr_refclk";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .gpon_lck2ref_control = "gpon_lck2ref_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .iqclk_mux_sel = "power_down";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .is_cascaded_pll = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lck2ref_delay_control = "lck2ref_delay_2";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lf_resistor_pd = "lf_pd_setting0";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lf_resistor_pfd = "lf_pfd_setting2";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lf_ripple_cap = "lf_no_ripple";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .loop_filter_bias_select = "lpflt_bias_7";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .loopback_mode = "loopback_disabled";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lpd_counter = 5'b01000;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .lpfd_counter = 5'b00001;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .ltd_ltr_micro_controller_select = "ltd_ltr_pcs";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .m_counter = 40;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .n_counter = 1;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .n_counter_scratch = 6'b000001;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .optimal = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .output_clock_frequency = "625000000 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pcie_gen = "non_pcie";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pd_fastlock_mode = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pd_l_counter = 8;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pfd_l_counter = 1;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pm_speed_grade = "e2";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .pma_width = 10;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .position = "position_unknown";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .power_mode = "low_power";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .primary_use = "cdr";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .reference_clock_frequency = "125000000 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .requires_gt_capable_channel = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .reverse_serial_loopback = "no_loopback";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_input_freq_range = 8'b00000000;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_v2i_enable = "true";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_vco_reset = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_vco_speed = 5'b00011;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_vco_speed_fix = 8'b00111100;
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .set_cdr_vco_speed_pciegen3 = "cdr_vco_max_speedbin_pciegen3";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .side = "side_unknown";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .sup_mode = "user_mode";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .top_or_bottom = "tb_unknown";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .tx_pll_prot_mode = "txpll_unused";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .txpll_hclk_driver_enable = "false";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .uc_cru_rstb = "cdr_lf_reset_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .uc_ro_cal = "uc_ro_cal_on";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .uc_ro_cal_status = "uc_ro_cal_notdone";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .vco_freq = "5000000000 hz";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .vco_overrange_voltage = "vco_overrange_off";
defparam \gen_twentynm_hssi_pma_channel_pll.inst_twentynm_hssi_pma_channel_pll .vco_underrange_voltage = "vco_underange_off";

twentynm_hssi_pma_cdr_refclk_select_mux \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux (
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.core_refclk(gnd),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.iqtxrxclk({gnd,gnd,gnd,gnd,gnd,gnd}),
	.ref_iqclk({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,in_ref_iqclk[0]}),
	.blockselect(out_blockselect_pma_cdr_refclk),
	.refclk(w_pma_cdr_refclk_refclk),
	.rx_det_clk(w_pma_cdr_refclk_rx_det_clk),
	.avmmreaddata(\gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux_AVMMREADDATA_bus ));
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .cdr_clkin_scratch0_src = "cdr_clkin_scratch0_src_refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .cdr_clkin_scratch1_src = "cdr_clkin_scratch1_src_refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .cdr_clkin_scratch2_src = "cdr_clkin_scratch2_src_refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .cdr_clkin_scratch3_src = "cdr_clkin_scratch3_src_refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .cdr_clkin_scratch4_src = "cdr_clkin_scratch4_src_refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .inclk0_logical_to_physical_mapping = "ref_iqclk0";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .inclk1_logical_to_physical_mapping = "power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .inclk2_logical_to_physical_mapping = "power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .inclk3_logical_to_physical_mapping = "power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .inclk4_logical_to_physical_mapping = "power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .powerdown_mode = "powerup";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .receiver_detect_src = "iqclk_src";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .refclk_select = "ref_iqclk0";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xmux_refclk_src = "refclk_iqclk";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_iqclk_sel = "power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_scratch0_src = "scratch0_power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_scratch1_src = "scratch1_power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_scratch2_src = "scratch2_power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_scratch3_src = "scratch3_power_down";
defparam \gen_twentynm_hssi_pma_cdr_refclk_select_mux.inst_twentynm_hssi_pma_cdr_refclk_select_mux .xpm_iqref_mux_scratch4_src = "scratch4_power_down";

twentynm_hssi_pma_adaptation \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation (
	.adapt_reset(gnd),
	.adapt_start(gnd),
	.avmmclk(in_avmmclk),
	.avmmread(in_avmmread),
	.avmmrstn(in_avmmrstn),
	.avmmwrite(in_avmmwrite),
	.deser_clk(w_pma_rx_deser_adapt_clk),
	.deser_odi_clk(gnd),
	.global_pipe_se(vcc),
	.radp_ctle_hold_en(),
	.radp_ctle_patt_en(),
	.radp_ctle_preset_sel(),
	.radp_enable_max_lfeq_scale(),
	.radp_lfeq_hold_en(),
	.radp_vga_polarity(),
	.rx_pllfreqlock(out_rxpll_lock),
	.scan_clk(gnd),
	.test_mode(vcc),
	.test_se(vcc),
	.avmmaddress({in_avmmaddress[8],in_avmmaddress[7],in_avmmaddress[6],in_avmmaddress[5],in_avmmaddress[4],in_avmmaddress[3],in_avmmaddress[2],in_avmmaddress[1],in_avmmaddress[0]}),
	.avmmwritedata({in_avmmwritedata[7],in_avmmwritedata[6],in_avmmwritedata[5],in_avmmwritedata[4],in_avmmwritedata[3],in_avmmwritedata[2],in_avmmwritedata[1],in_avmmwritedata[0]}),
	.deser_data({\w_pma_rx_deser_data[63] ,\w_pma_rx_deser_data[62] ,\w_pma_rx_deser_data[61] ,\w_pma_rx_deser_data[60] ,\w_pma_rx_deser_data[59] ,\w_pma_rx_deser_data[58] ,\w_pma_rx_deser_data[57] ,\w_pma_rx_deser_data[56] ,\w_pma_rx_deser_data[55] ,\w_pma_rx_deser_data[54] ,
\w_pma_rx_deser_data[53] ,\w_pma_rx_deser_data[52] ,\w_pma_rx_deser_data[51] ,\w_pma_rx_deser_data[50] ,\w_pma_rx_deser_data[49] ,\w_pma_rx_deser_data[48] ,\w_pma_rx_deser_data[47] ,\w_pma_rx_deser_data[46] ,\w_pma_rx_deser_data[45] ,\w_pma_rx_deser_data[44] ,
\w_pma_rx_deser_data[43] ,\w_pma_rx_deser_data[42] ,\w_pma_rx_deser_data[41] ,\w_pma_rx_deser_data[40] ,\w_pma_rx_deser_data[39] ,\w_pma_rx_deser_data[38] ,\w_pma_rx_deser_data[37] ,\w_pma_rx_deser_data[36] ,\w_pma_rx_deser_data[35] ,\w_pma_rx_deser_data[34] ,
\w_pma_rx_deser_data[33] ,\w_pma_rx_deser_data[32] ,\w_pma_rx_deser_data[31] ,\w_pma_rx_deser_data[30] ,\w_pma_rx_deser_data[29] ,\w_pma_rx_deser_data[28] ,\w_pma_rx_deser_data[27] ,\w_pma_rx_deser_data[26] ,\w_pma_rx_deser_data[25] ,\w_pma_rx_deser_data[24] ,
\w_pma_rx_deser_data[23] ,\w_pma_rx_deser_data[22] ,\w_pma_rx_deser_data[21] ,\w_pma_rx_deser_data[20] ,\w_pma_rx_deser_data[19] ,\w_pma_rx_deser_data[18] ,\w_pma_rx_deser_data[17] ,\w_pma_rx_deser_data[16] ,\w_pma_rx_deser_data[15] ,\w_pma_rx_deser_data[14] ,
\w_pma_rx_deser_data[13] ,\w_pma_rx_deser_data[12] ,\w_pma_rx_deser_data[11] ,\w_pma_rx_deser_data[10] ,\w_pma_rx_deser_data[9] ,\w_pma_rx_deser_data[8] ,\w_pma_rx_deser_data[7] ,\w_pma_rx_deser_data[6] ,\w_pma_rx_deser_data[5] ,\w_pma_rx_deser_data[4] ,
\w_pma_rx_deser_data[3] ,\w_pma_rx_deser_data[2] ,\w_pma_rx_deser_data[1] ,\w_pma_rx_deser_data[0] }),
	.deser_error({\w_pma_rx_deser_error_deser[63] ,\w_pma_rx_deser_error_deser[62] ,\w_pma_rx_deser_error_deser[61] ,\w_pma_rx_deser_error_deser[60] ,\w_pma_rx_deser_error_deser[59] ,\w_pma_rx_deser_error_deser[58] ,\w_pma_rx_deser_error_deser[57] ,\w_pma_rx_deser_error_deser[56] ,
\w_pma_rx_deser_error_deser[55] ,\w_pma_rx_deser_error_deser[54] ,\w_pma_rx_deser_error_deser[53] ,\w_pma_rx_deser_error_deser[52] ,\w_pma_rx_deser_error_deser[51] ,\w_pma_rx_deser_error_deser[50] ,\w_pma_rx_deser_error_deser[49] ,\w_pma_rx_deser_error_deser[48] ,
\w_pma_rx_deser_error_deser[47] ,\w_pma_rx_deser_error_deser[46] ,\w_pma_rx_deser_error_deser[45] ,\w_pma_rx_deser_error_deser[44] ,\w_pma_rx_deser_error_deser[43] ,\w_pma_rx_deser_error_deser[42] ,\w_pma_rx_deser_error_deser[41] ,\w_pma_rx_deser_error_deser[40] ,
\w_pma_rx_deser_error_deser[39] ,\w_pma_rx_deser_error_deser[38] ,\w_pma_rx_deser_error_deser[37] ,\w_pma_rx_deser_error_deser[36] ,\w_pma_rx_deser_error_deser[35] ,\w_pma_rx_deser_error_deser[34] ,\w_pma_rx_deser_error_deser[33] ,\w_pma_rx_deser_error_deser[32] ,
\w_pma_rx_deser_error_deser[31] ,\w_pma_rx_deser_error_deser[30] ,\w_pma_rx_deser_error_deser[29] ,\w_pma_rx_deser_error_deser[28] ,\w_pma_rx_deser_error_deser[27] ,\w_pma_rx_deser_error_deser[26] ,\w_pma_rx_deser_error_deser[25] ,\w_pma_rx_deser_error_deser[24] ,
\w_pma_rx_deser_error_deser[23] ,\w_pma_rx_deser_error_deser[22] ,\w_pma_rx_deser_error_deser[21] ,\w_pma_rx_deser_error_deser[20] ,\w_pma_rx_deser_error_deser[19] ,\w_pma_rx_deser_error_deser[18] ,\w_pma_rx_deser_error_deser[17] ,\w_pma_rx_deser_error_deser[16] ,
\w_pma_rx_deser_error_deser[15] ,\w_pma_rx_deser_error_deser[14] ,\w_pma_rx_deser_error_deser[13] ,\w_pma_rx_deser_error_deser[12] ,\w_pma_rx_deser_error_deser[11] ,\w_pma_rx_deser_error_deser[10] ,\w_pma_rx_deser_error_deser[9] ,\w_pma_rx_deser_error_deser[8] ,
\w_pma_rx_deser_error_deser[7] ,\w_pma_rx_deser_error_deser[6] ,\w_pma_rx_deser_error_deser[5] ,\w_pma_rx_deser_error_deser[4] ,\w_pma_rx_deser_error_deser[3] ,\w_pma_rx_deser_error_deser[2] ,\w_pma_rx_deser_error_deser[1] ,\w_pma_rx_deser_error_deser[0] }),
	.deser_odi({\w_pma_rx_deser_odi_dout[63] ,\w_pma_rx_deser_odi_dout[62] ,\w_pma_rx_deser_odi_dout[61] ,\w_pma_rx_deser_odi_dout[60] ,\w_pma_rx_deser_odi_dout[59] ,\w_pma_rx_deser_odi_dout[58] ,\w_pma_rx_deser_odi_dout[57] ,\w_pma_rx_deser_odi_dout[56] ,
\w_pma_rx_deser_odi_dout[55] ,\w_pma_rx_deser_odi_dout[54] ,\w_pma_rx_deser_odi_dout[53] ,\w_pma_rx_deser_odi_dout[52] ,\w_pma_rx_deser_odi_dout[51] ,\w_pma_rx_deser_odi_dout[50] ,\w_pma_rx_deser_odi_dout[49] ,\w_pma_rx_deser_odi_dout[48] ,
\w_pma_rx_deser_odi_dout[47] ,\w_pma_rx_deser_odi_dout[46] ,\w_pma_rx_deser_odi_dout[45] ,\w_pma_rx_deser_odi_dout[44] ,\w_pma_rx_deser_odi_dout[43] ,\w_pma_rx_deser_odi_dout[42] ,\w_pma_rx_deser_odi_dout[41] ,\w_pma_rx_deser_odi_dout[40] ,
\w_pma_rx_deser_odi_dout[39] ,\w_pma_rx_deser_odi_dout[38] ,\w_pma_rx_deser_odi_dout[37] ,\w_pma_rx_deser_odi_dout[36] ,\w_pma_rx_deser_odi_dout[35] ,\w_pma_rx_deser_odi_dout[34] ,\w_pma_rx_deser_odi_dout[33] ,\w_pma_rx_deser_odi_dout[32] ,
\w_pma_rx_deser_odi_dout[31] ,\w_pma_rx_deser_odi_dout[30] ,\w_pma_rx_deser_odi_dout[29] ,\w_pma_rx_deser_odi_dout[28] ,\w_pma_rx_deser_odi_dout[27] ,\w_pma_rx_deser_odi_dout[26] ,\w_pma_rx_deser_odi_dout[25] ,\w_pma_rx_deser_odi_dout[24] ,
\w_pma_rx_deser_odi_dout[23] ,\w_pma_rx_deser_odi_dout[22] ,\w_pma_rx_deser_odi_dout[21] ,\w_pma_rx_deser_odi_dout[20] ,\w_pma_rx_deser_odi_dout[19] ,\w_pma_rx_deser_odi_dout[18] ,\w_pma_rx_deser_odi_dout[17] ,\w_pma_rx_deser_odi_dout[16] ,
\w_pma_rx_deser_odi_dout[15] ,\w_pma_rx_deser_odi_dout[14] ,\w_pma_rx_deser_odi_dout[13] ,\w_pma_rx_deser_odi_dout[12] ,\w_pma_rx_deser_odi_dout[11] ,\w_pma_rx_deser_odi_dout[10] ,\w_pma_rx_deser_odi_dout[9] ,\w_pma_rx_deser_odi_dout[8] ,
\w_pma_rx_deser_odi_dout[7] ,\w_pma_rx_deser_odi_dout[6] ,\w_pma_rx_deser_odi_dout[5] ,\w_pma_rx_deser_odi_dout[4] ,\w_pma_rx_deser_odi_dout[3] ,\w_pma_rx_deser_odi_dout[2] ,\w_pma_rx_deser_odi_dout[1] ,\w_pma_rx_deser_odi_dout[0] }),
	.i_rxpreset({gnd,gnd,gnd}),
	.scan_in({gnd,gnd,gnd,vcc,in_eye_monitor[5],in_eye_monitor[4],in_eye_monitor[3],in_eye_monitor[2],in_eye_monitor[1],in_eye_monitor[0]}),
	.blockselect(out_blockselect_pma_adapt),
	.dfe_adapt_en(w_pma_adapt_dfe_adapt_en),
	.dfe_adp_clk(w_pma_adapt_dfe_adp_clk),
	.dfe_fltap1_sgn(w_pma_adapt_dfe_fltap1_sgn),
	.dfe_fltap2_sgn(w_pma_adapt_dfe_fltap2_sgn),
	.dfe_fltap3_sgn(w_pma_adapt_dfe_fltap3_sgn),
	.dfe_fltap4_sgn(w_pma_adapt_dfe_fltap4_sgn),
	.dfe_fltap_bypdeser(w_pma_adapt_dfe_fltap_bypdeser),
	.dfe_fxtap2_sgn(w_pma_adapt_dfe_fxtap2_sgn),
	.dfe_fxtap3_sgn(w_pma_adapt_dfe_fxtap3_sgn),
	.dfe_fxtap4_sgn(w_pma_adapt_dfe_fxtap4_sgn),
	.dfe_fxtap5_sgn(w_pma_adapt_dfe_fxtap5_sgn),
	.dfe_fxtap6_sgn(w_pma_adapt_dfe_fxtap6_sgn),
	.dfe_fxtap7_sgn(w_pma_adapt_dfe_fxtap7_sgn),
	.dfe_spec_disable(w_pma_adapt_dfe_spec_disable),
	.dfe_spec_sign_sel(w_pma_adapt_dfe_spec_sign_sel),
	.dfe_vref_sign_sel(w_pma_adapt_dfe_vref_sign_sel),
	.avmmreaddata(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_AVMMREADDATA_bus ),
	.ctle_acgain_4s(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_ACGAIN_4S_bus ),
	.ctle_eqz_1s_sel(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_EQZ_1S_SEL_bus ),
	.ctle_lfeq_fb_sel(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_CTLE_LFEQ_FB_SEL_bus ),
	.dfe_fltap1(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP1_bus ),
	.dfe_fltap2(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP2_bus ),
	.dfe_fltap3(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP3_bus ),
	.dfe_fltap4(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP4_bus ),
	.dfe_fltap_position(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FLTAP_POSITION_bus ),
	.dfe_fxtap1(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP1_bus ),
	.dfe_fxtap2(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP2_bus ),
	.dfe_fxtap3(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP3_bus ),
	.dfe_fxtap4(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP4_bus ),
	.dfe_fxtap5(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP5_bus ),
	.dfe_fxtap6(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP6_bus ),
	.dfe_fxtap7(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_DFE_FXTAP7_bus ),
	.odi_vref(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_ODI_VREF_bus ),
	.scan_out(),
	.status_bus(),
	.vga_sel(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VGA_SEL_bus ),
	.vref_sel(\gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation_VREF_SEL_bus ));
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adapt_dfe_control_sel = "r_adapt_dfe_control_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adapt_dfe_sel = "r_adapt_dfe_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adapt_mode = "manual";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adapt_vga_sel = "r_adapt_vga_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adapt_vref_sel = "r_adapt_vref_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_1s_ctle_bypass = "radp_1s_ctle_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_4s_ctle_bypass = "radp_4s_ctle_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_adapt_control_sel = "radp_adapt_control_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_adapt_rstn = "radp_adapt_rstn_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_adapt_start = "radp_adapt_start_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_auxpath_en = "radp_bist_auxpath_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_count_rstn = "radp_bist_count_rstn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_datapath_en = "radp_bist_datapath_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_mode = "radp_bist_mode_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_odi_dfe_sel = "radp_bist_odi_dfe_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_bist_spec_en = "radp_bist_spec_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_control_mux_bypass = "radp_control_mux_bypass_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_acgain_4s = "radp_ctle_acgain_4s_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_adapt_bw = "radp_ctle_adapt_bw_3";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_adapt_cycle_window = "radp_ctle_adapt_cycle_window_7";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_adapt_oneshot = "radp_ctle_adapt_oneshot_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_en = "radp_ctle_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_eqz_1s_sel = "radp_ctle_eqz_1s_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_force_spec_sign = "radp_ctle_force_spec_sign_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_hold_en = "radp_ctle_not_held";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_load = "radp_ctle_load_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_load_value = "radp_ctle_load_value_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_scale = "radp_ctle_scale_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_scale_en = "radp_ctle_scale_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_spec_sign = "radp_ctle_spec_sign_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_sweep_direction = "radp_ctle_sweep_direction_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_threshold = "radp_ctle_threshold_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_threshold_en = "radp_ctle_threshold_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_vref_polarity = "radp_ctle_vref_polarity_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_ctle_window = "radp_ctle_window_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_bw = "radp_dfe_bw_3";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_clkout_div_sel = "radp_dfe_clkout_div_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_cycle = "radp_dfe_cycle_6";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fltap_bypass = "radp_dfe_fltap_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fltap_en = "radp_dfe_fltap_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fltap_hold_en = "radp_dfe_fltap_not_held";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fltap_load = "radp_dfe_fltap_load_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fltap_position = "radp_dfe_fltap_position_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_force_spec_sign = "radp_dfe_force_spec_sign_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap1 = "radp_dfe_fxtap1_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap10 = "radp_dfe_fxtap10_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap10_sgn = "radp_dfe_fxtap10_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap11 = "radp_dfe_fxtap11_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap11_sgn = "radp_dfe_fxtap11_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap2 = "radp_dfe_fxtap2_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap2_sgn = "radp_dfe_fxtap2_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap3 = "radp_dfe_fxtap3_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap3_sgn = "radp_dfe_fxtap3_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap4 = "radp_dfe_fxtap4_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap4_sgn = "radp_dfe_fxtap4_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap5 = "radp_dfe_fxtap5_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap5_sgn = "radp_dfe_fxtap5_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap6 = "radp_dfe_fxtap6_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap6_sgn = "radp_dfe_fxtap6_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap7 = "radp_dfe_fxtap7_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap7_sgn = "radp_dfe_fxtap7_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap8 = "radp_dfe_fxtap8_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap8_sgn = "radp_dfe_fxtap8_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap9 = "radp_dfe_fxtap9_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap9_sgn = "radp_dfe_fxtap9_sgn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap_bypass = "radp_dfe_fxtap_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap_en = "radp_dfe_fxtap_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap_hold_en = "radp_dfe_fxtap_not_held";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_fxtap_load = "radp_dfe_fxtap_load_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_mode = "radp_dfe_mode_4";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_spec_sign = "radp_dfe_spec_sign_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_dfe_vref_polarity = "radp_dfe_vref_polarity_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_force_freqlock = "radp_force_freqlock_off";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_frame_capture = "radp_frame_capture_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_frame_en = "radp_frame_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_frame_odi_sel = "radp_frame_odi_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_frame_out_sel = "radp_frame_out_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_lfeq_fb_sel = "radp_lfeq_fb_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_mode = "radp_mode_8";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_odi_control_sel = "radp_odi_control_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_onetime_dfe = "radp_onetime_dfe_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_spec_avg_window = "radp_spec_avg_window_4";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_spec_trans_filter = "radp_spec_trans_filter_2";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_status_sel = "radp_status_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_bypass = "radp_vga_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_en = "radp_vga_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_load = "radp_vga_load_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_polarity = "radp_vga_polarity_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_sel = "radp_vga_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_sweep_direction = "radp_vga_sweep_direction_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vga_threshold = "radp_vga_threshold_4";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_bw = "radp_vref_bw_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_bypass = "radp_vref_bypass_1";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_cycle = "radp_vref_cycle_6";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_dfe_spec_en = "radp_vref_dfe_spec_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_en = "radp_vref_disable";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_hold_en = "radp_vref_not_held";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_load = "radp_vref_load_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_polarity = "radp_vref_polarity_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_sel = "radp_vref_sel_21";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .adp_vref_vga_level = "radp_vref_vga_level_13";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .datarate = "1250000000 bps";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .initial_settings = "true";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_count_threshold = "rodi_count_threshold_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_dfe_spec_en = "rodi_dfe_spec_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_en = "rodi_en_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_mode = "rodi_mode_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_rstn = "rodi_rstn_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_spec_sel = "rodi_spec_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_start = "rodi_start_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .odi_vref_sel = "rodi_vref_sel_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .optimal = "false";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .prot_mode = "basic_rx";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .rrx_pcie_eqz = "rrx_pcie_eqz_0";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .silicon_rev = "20nm5";
defparam \gen_twentynm_hssi_pma_adaptation.inst_twentynm_hssi_pma_adaptation .sup_mode = "user_mode";

endmodule

module wr_arria10_e3p1_det_phy_twentynm_xcvr_avmm (
	pcs_blockselect_rx_pcs_pld_if,
	pcs_avmmreaddata_rx_pcs_pld_if,
	chnl_pll_avmm_clk,
	pld_cal_done,
	chnl_pll_avmm_read,
	chnl_pll_avmm_rstn,
	chnl_pll_avmm_write,
	avmm_readdata,
	chnl_pll_avmm_address,
	chnl_pll_avmm_writedata,
	pcs_blockselect_com_pcs_pld_if,
	pcs_avmmreaddata_com_pcs_pld_if,
	pcs_blockselect_tx_pcs_pld_if,
	pcs_avmmreaddata_tx_pcs_pld_if,
	pma_blockselect_tx_buf,
	pma_avmmreaddata_tx_buf,
	pcs_blockselect_10g_rx_pcs,
	pcs_avmmreaddata_10g_rx_pcs,
	pcs_blockselect_8g_rx_pcs,
	pcs_avmmreaddata_8g_rx_pcs,
	pcs_blockselect_pipe_gen1_2,
	pcs_avmmreaddata_pipe_gen1_2,
	pcs_blockselect_krfec_rx_pcs,
	pcs_avmmreaddata_krfec_rx_pcs,
	pcs_blockselect_rx_pcs_pma_if,
	pcs_avmmreaddata_rx_pcs_pma_if,
	pma_blockselect_tx_ser,
	pma_avmmreaddata_tx_ser,
	pma_blockselect_tx_cgb,
	pma_avmmreaddata_tx_cgb,
	pma_blockselect_rx_deser,
	pma_avmmreaddata_rx_deser,
	pma_blockselect_rx_buf,
	pma_avmmreaddata_rx_buf,
	pma_blockselect_rx_sd,
	pma_avmmreaddata_rx_sd,
	pma_blockselect_rx_odi,
	pma_avmmreaddata_rx_odi,
	pma_blockselect_rx_dfe,
	pma_avmmreaddata_rx_dfe,
	pma_blockselect_cdr_pll,
	pma_avmmreaddata_cdr_pll,
	pma_blockselect_cdr_refclk_select,
	pma_avmmreaddata_cdr_refclk_select,
	pma_blockselect_pma_adapt,
	pma_avmmreaddata_pma_adapt,
	pcs_blockselect_8g_tx_pcs,
	pcs_avmmreaddata_8g_tx_pcs,
	pcs_blockselect_10g_tx_pcs,
	pcs_avmmreaddata_10g_tx_pcs,
	pcs_blockselect_gen3_rx_pcs,
	pcs_avmmreaddata_gen3_rx_pcs,
	pcs_blockselect_pipe_gen3,
	pcs_avmmreaddata_pipe_gen3,
	pcs_blockselect_gen3_tx_pcs,
	pcs_avmmreaddata_gen3_tx_pcs,
	pcs_blockselect_krfec_tx_pcs,
	pcs_avmmreaddata_krfec_tx_pcs,
	pcs_blockselect_fifo_rx_pcs,
	pcs_avmmreaddata_fifo_rx_pcs,
	pcs_blockselect_fifo_tx_pcs,
	pcs_avmmreaddata_fifo_tx_pcs,
	pcs_blockselect_com_pcs_pma_if,
	pcs_avmmreaddata_com_pcs_pma_if,
	pcs_blockselect_tx_pcs_pma_if,
	pcs_avmmreaddata_tx_pcs_pma_if,
	avmm_waitrequest_0,
	avmm_read,
	reconfig_clk_0,
	avmm_write,
	avmm_address,
	avmm_writedata,
	reconfig_reset_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] pcs_blockselect_rx_pcs_pld_if;
input 	[7:0] pcs_avmmreaddata_rx_pcs_pld_if;
output 	[0:0] chnl_pll_avmm_clk;
output 	[0:0] pld_cal_done;
output 	[0:0] chnl_pll_avmm_read;
output 	[0:0] chnl_pll_avmm_rstn;
output 	[0:0] chnl_pll_avmm_write;
output 	[7:0] avmm_readdata;
output 	[8:0] chnl_pll_avmm_address;
output 	[7:0] chnl_pll_avmm_writedata;
input 	[0:0] pcs_blockselect_com_pcs_pld_if;
input 	[7:0] pcs_avmmreaddata_com_pcs_pld_if;
input 	[0:0] pcs_blockselect_tx_pcs_pld_if;
input 	[7:0] pcs_avmmreaddata_tx_pcs_pld_if;
input 	[0:0] pma_blockselect_tx_buf;
input 	[7:0] pma_avmmreaddata_tx_buf;
input 	[0:0] pcs_blockselect_10g_rx_pcs;
input 	[7:0] pcs_avmmreaddata_10g_rx_pcs;
input 	[0:0] pcs_blockselect_8g_rx_pcs;
input 	[7:0] pcs_avmmreaddata_8g_rx_pcs;
input 	[0:0] pcs_blockselect_pipe_gen1_2;
input 	[7:0] pcs_avmmreaddata_pipe_gen1_2;
input 	[0:0] pcs_blockselect_krfec_rx_pcs;
input 	[7:0] pcs_avmmreaddata_krfec_rx_pcs;
input 	[0:0] pcs_blockselect_rx_pcs_pma_if;
input 	[7:0] pcs_avmmreaddata_rx_pcs_pma_if;
input 	[0:0] pma_blockselect_tx_ser;
input 	[7:0] pma_avmmreaddata_tx_ser;
input 	[0:0] pma_blockselect_tx_cgb;
input 	[7:0] pma_avmmreaddata_tx_cgb;
input 	[0:0] pma_blockselect_rx_deser;
input 	[7:0] pma_avmmreaddata_rx_deser;
input 	[0:0] pma_blockselect_rx_buf;
input 	[7:0] pma_avmmreaddata_rx_buf;
input 	[0:0] pma_blockselect_rx_sd;
input 	[7:0] pma_avmmreaddata_rx_sd;
input 	[0:0] pma_blockselect_rx_odi;
input 	[7:0] pma_avmmreaddata_rx_odi;
input 	[0:0] pma_blockselect_rx_dfe;
input 	[7:0] pma_avmmreaddata_rx_dfe;
input 	[0:0] pma_blockselect_cdr_pll;
input 	[7:0] pma_avmmreaddata_cdr_pll;
input 	[0:0] pma_blockselect_cdr_refclk_select;
input 	[7:0] pma_avmmreaddata_cdr_refclk_select;
input 	[0:0] pma_blockselect_pma_adapt;
input 	[7:0] pma_avmmreaddata_pma_adapt;
input 	[0:0] pcs_blockselect_8g_tx_pcs;
input 	[7:0] pcs_avmmreaddata_8g_tx_pcs;
input 	[0:0] pcs_blockselect_10g_tx_pcs;
input 	[7:0] pcs_avmmreaddata_10g_tx_pcs;
input 	[0:0] pcs_blockselect_gen3_rx_pcs;
input 	[7:0] pcs_avmmreaddata_gen3_rx_pcs;
input 	[0:0] pcs_blockselect_pipe_gen3;
input 	[7:0] pcs_avmmreaddata_pipe_gen3;
input 	[0:0] pcs_blockselect_gen3_tx_pcs;
input 	[7:0] pcs_avmmreaddata_gen3_tx_pcs;
input 	[0:0] pcs_blockselect_krfec_tx_pcs;
input 	[7:0] pcs_avmmreaddata_krfec_tx_pcs;
input 	[0:0] pcs_blockselect_fifo_rx_pcs;
input 	[7:0] pcs_avmmreaddata_fifo_rx_pcs;
input 	[0:0] pcs_blockselect_fifo_tx_pcs;
input 	[7:0] pcs_avmmreaddata_fifo_tx_pcs;
input 	[0:0] pcs_blockselect_com_pcs_pma_if;
input 	[7:0] pcs_avmmreaddata_com_pcs_pma_if;
input 	[0:0] pcs_blockselect_tx_pcs_pma_if;
input 	[7:0] pcs_avmmreaddata_tx_pcs_pma_if;
output 	avmm_waitrequest_0;
input 	[0:0] avmm_read;
input 	reconfig_clk_0;
input 	[0:0] avmm_write;
input 	[8:0] avmm_address;
input 	[7:0] avmm_writedata;
input 	reconfig_reset_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ;
wire \avmm_busy[0] ;
wire \avmm_busy_r1[0]~q ;
wire \avmm_busy_r2[0]~q ;
wire \avmm_waitrequest_write_int~0_combout ;
wire \avmm_waitrequest_write_int~1_combout ;
wire \avmm_waitrequest_write_int~2_combout ;
wire \avmm_waitrequest_write_int[0]~q ;
wire \avmm_read_r[0]~q ;
wire \avmm_read_cycles_cnt~2_combout ;
wire \avmm_read_cycles_cnt[0]~q ;
wire \avmm_read_cycles_cnt~1_combout ;
wire \avmm_read_cycles_cnt[2]~q ;
wire \avmm_read_cycles_cnt~0_combout ;
wire \avmm_read_cycles_cnt[1]~q ;

wire [7:0] \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus ;
wire [8:0] \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus ;
wire [7:0] \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus ;

assign chnl_pll_avmm_writedata[0] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [0];
assign chnl_pll_avmm_writedata[1] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [1];
assign chnl_pll_avmm_writedata[2] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [2];
assign chnl_pll_avmm_writedata[3] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [3];
assign chnl_pll_avmm_writedata[4] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [4];
assign chnl_pll_avmm_writedata[5] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [5];
assign chnl_pll_avmm_writedata[6] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [6];
assign chnl_pll_avmm_writedata[7] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus [7];

assign chnl_pll_avmm_address[0] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [0];
assign chnl_pll_avmm_address[1] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [1];
assign chnl_pll_avmm_address[2] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [2];
assign chnl_pll_avmm_address[3] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [3];
assign chnl_pll_avmm_address[4] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [4];
assign chnl_pll_avmm_address[5] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [5];
assign chnl_pll_avmm_address[6] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [6];
assign chnl_pll_avmm_address[7] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [7];
assign chnl_pll_avmm_address[8] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus [8];

assign avmm_readdata[0] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [0];
assign avmm_readdata[1] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [1];
assign avmm_readdata[2] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [2];
assign avmm_readdata[3] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [3];
assign avmm_readdata[4] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [4];
assign avmm_readdata[5] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [5];
assign avmm_readdata[6] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [6];
assign avmm_readdata[7] = \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus [7];

wr_arria10_e3p1_det_phy_alt_xcvr_resync \avmm_atom_insts[0].avmm_reset_sync_inst (
	.resync_chains0sync_r_1(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.clk(reconfig_clk_0),
	.reconfig_reset_0(reconfig_reset_0));

twentynm_hssi_avmm_if \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst (
	.avmmclk(reconfig_clk_0),
	.avmmread(avmm_read[0]),
	.avmmrequest(vcc),
	.avmmreservedin(),
	.avmmrstn(vcc),
	.avmmwrite(avmm_write[0]),
	.scanmoden(vcc),
	.scanshiftn(vcc),
	.avmmaddress({avmm_address[8],avmm_address[7],avmm_address[6],avmm_address[5],avmm_address[4],avmm_address[3],avmm_address[2],avmm_address[1],avmm_address[0]}),
	.avmmwritedata({avmm_writedata[7],avmm_writedata[6],avmm_writedata[5],avmm_writedata[4],avmm_writedata[3],avmm_writedata[2],avmm_writedata[1],avmm_writedata[0]}),
	.blockselect({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,pcs_blockselect_tx_pcs_pma_if[0],pcs_blockselect_com_pcs_pma_if[0],pcs_blockselect_rx_pcs_pma_if[0],pcs_blockselect_tx_pcs_pld_if[0],pcs_blockselect_com_pcs_pld_if[0],
pcs_blockselect_rx_pcs_pld_if[0],pcs_blockselect_fifo_tx_pcs[0],pcs_blockselect_fifo_rx_pcs[0],pcs_blockselect_krfec_tx_pcs[0],pcs_blockselect_krfec_rx_pcs[0],pcs_blockselect_gen3_tx_pcs[0],pcs_blockselect_pipe_gen3[0],pcs_blockselect_gen3_rx_pcs[0],pcs_blockselect_10g_tx_pcs[0],
pcs_blockselect_10g_rx_pcs[0],pcs_blockselect_8g_tx_pcs[0],pcs_blockselect_pipe_gen1_2[0],pcs_blockselect_8g_rx_pcs[0],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,pma_blockselect_pma_adapt[0],pma_blockselect_cdr_refclk_select[0],pma_blockselect_cdr_pll[0],pma_blockselect_rx_dfe[0],pma_blockselect_rx_odi[0],
pma_blockselect_rx_sd[0],pma_blockselect_rx_buf[0],pma_blockselect_rx_deser[0],pma_blockselect_tx_buf[0],pma_blockselect_tx_cgb[0],pma_blockselect_tx_ser[0]}),
	.readdatachnl({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,pcs_avmmreaddata_tx_pcs_pma_if[7],pcs_avmmreaddata_tx_pcs_pma_if[6],pcs_avmmreaddata_tx_pcs_pma_if[5],pcs_avmmreaddata_tx_pcs_pma_if[4],pcs_avmmreaddata_tx_pcs_pma_if[3],pcs_avmmreaddata_tx_pcs_pma_if[2],pcs_avmmreaddata_tx_pcs_pma_if[1],pcs_avmmreaddata_tx_pcs_pma_if[0],
pcs_avmmreaddata_com_pcs_pma_if[7],pcs_avmmreaddata_com_pcs_pma_if[6],pcs_avmmreaddata_com_pcs_pma_if[5],pcs_avmmreaddata_com_pcs_pma_if[4],pcs_avmmreaddata_com_pcs_pma_if[3],pcs_avmmreaddata_com_pcs_pma_if[2],pcs_avmmreaddata_com_pcs_pma_if[1],pcs_avmmreaddata_com_pcs_pma_if[0],
pcs_avmmreaddata_rx_pcs_pma_if[7],pcs_avmmreaddata_rx_pcs_pma_if[6],pcs_avmmreaddata_rx_pcs_pma_if[5],pcs_avmmreaddata_rx_pcs_pma_if[4],pcs_avmmreaddata_rx_pcs_pma_if[3],pcs_avmmreaddata_rx_pcs_pma_if[2],pcs_avmmreaddata_rx_pcs_pma_if[1],pcs_avmmreaddata_rx_pcs_pma_if[0],
pcs_avmmreaddata_tx_pcs_pld_if[7],pcs_avmmreaddata_tx_pcs_pld_if[6],pcs_avmmreaddata_tx_pcs_pld_if[5],pcs_avmmreaddata_tx_pcs_pld_if[4],pcs_avmmreaddata_tx_pcs_pld_if[3],pcs_avmmreaddata_tx_pcs_pld_if[2],pcs_avmmreaddata_tx_pcs_pld_if[1],pcs_avmmreaddata_tx_pcs_pld_if[0],
pcs_avmmreaddata_com_pcs_pld_if[7],pcs_avmmreaddata_com_pcs_pld_if[6],pcs_avmmreaddata_com_pcs_pld_if[5],pcs_avmmreaddata_com_pcs_pld_if[4],pcs_avmmreaddata_com_pcs_pld_if[3],pcs_avmmreaddata_com_pcs_pld_if[2],pcs_avmmreaddata_com_pcs_pld_if[1],pcs_avmmreaddata_com_pcs_pld_if[0],
pcs_avmmreaddata_rx_pcs_pld_if[7],pcs_avmmreaddata_rx_pcs_pld_if[6],pcs_avmmreaddata_rx_pcs_pld_if[5],pcs_avmmreaddata_rx_pcs_pld_if[4],pcs_avmmreaddata_rx_pcs_pld_if[3],pcs_avmmreaddata_rx_pcs_pld_if[2],pcs_avmmreaddata_rx_pcs_pld_if[1],pcs_avmmreaddata_rx_pcs_pld_if[0],
pcs_avmmreaddata_fifo_tx_pcs[7],pcs_avmmreaddata_fifo_tx_pcs[6],pcs_avmmreaddata_fifo_tx_pcs[5],pcs_avmmreaddata_fifo_tx_pcs[4],pcs_avmmreaddata_fifo_tx_pcs[3],pcs_avmmreaddata_fifo_tx_pcs[2],pcs_avmmreaddata_fifo_tx_pcs[1],pcs_avmmreaddata_fifo_tx_pcs[0],pcs_avmmreaddata_fifo_rx_pcs[7],
pcs_avmmreaddata_fifo_rx_pcs[6],pcs_avmmreaddata_fifo_rx_pcs[5],pcs_avmmreaddata_fifo_rx_pcs[4],pcs_avmmreaddata_fifo_rx_pcs[3],pcs_avmmreaddata_fifo_rx_pcs[2],pcs_avmmreaddata_fifo_rx_pcs[1],pcs_avmmreaddata_fifo_rx_pcs[0],pcs_avmmreaddata_krfec_tx_pcs[7],pcs_avmmreaddata_krfec_tx_pcs[6],
pcs_avmmreaddata_krfec_tx_pcs[5],pcs_avmmreaddata_krfec_tx_pcs[4],pcs_avmmreaddata_krfec_tx_pcs[3],pcs_avmmreaddata_krfec_tx_pcs[2],pcs_avmmreaddata_krfec_tx_pcs[1],pcs_avmmreaddata_krfec_tx_pcs[0],pcs_avmmreaddata_krfec_rx_pcs[7],pcs_avmmreaddata_krfec_rx_pcs[6],
pcs_avmmreaddata_krfec_rx_pcs[5],pcs_avmmreaddata_krfec_rx_pcs[4],pcs_avmmreaddata_krfec_rx_pcs[3],pcs_avmmreaddata_krfec_rx_pcs[2],pcs_avmmreaddata_krfec_rx_pcs[1],pcs_avmmreaddata_krfec_rx_pcs[0],pcs_avmmreaddata_gen3_tx_pcs[7],pcs_avmmreaddata_gen3_tx_pcs[6],
pcs_avmmreaddata_gen3_tx_pcs[5],pcs_avmmreaddata_gen3_tx_pcs[4],pcs_avmmreaddata_gen3_tx_pcs[3],pcs_avmmreaddata_gen3_tx_pcs[2],pcs_avmmreaddata_gen3_tx_pcs[1],pcs_avmmreaddata_gen3_tx_pcs[0],pcs_avmmreaddata_pipe_gen3[7],pcs_avmmreaddata_pipe_gen3[6],pcs_avmmreaddata_pipe_gen3[5],
pcs_avmmreaddata_pipe_gen3[4],pcs_avmmreaddata_pipe_gen3[3],pcs_avmmreaddata_pipe_gen3[2],pcs_avmmreaddata_pipe_gen3[1],pcs_avmmreaddata_pipe_gen3[0],pcs_avmmreaddata_gen3_rx_pcs[7],pcs_avmmreaddata_gen3_rx_pcs[6],pcs_avmmreaddata_gen3_rx_pcs[5],pcs_avmmreaddata_gen3_rx_pcs[4],
pcs_avmmreaddata_gen3_rx_pcs[3],pcs_avmmreaddata_gen3_rx_pcs[2],pcs_avmmreaddata_gen3_rx_pcs[1],pcs_avmmreaddata_gen3_rx_pcs[0],pcs_avmmreaddata_10g_tx_pcs[7],pcs_avmmreaddata_10g_tx_pcs[6],pcs_avmmreaddata_10g_tx_pcs[5],pcs_avmmreaddata_10g_tx_pcs[4],pcs_avmmreaddata_10g_tx_pcs[3],
pcs_avmmreaddata_10g_tx_pcs[2],pcs_avmmreaddata_10g_tx_pcs[1],pcs_avmmreaddata_10g_tx_pcs[0],pcs_avmmreaddata_10g_rx_pcs[7],pcs_avmmreaddata_10g_rx_pcs[6],pcs_avmmreaddata_10g_rx_pcs[5],pcs_avmmreaddata_10g_rx_pcs[4],pcs_avmmreaddata_10g_rx_pcs[3],pcs_avmmreaddata_10g_rx_pcs[2],
pcs_avmmreaddata_10g_rx_pcs[1],pcs_avmmreaddata_10g_rx_pcs[0],pcs_avmmreaddata_8g_tx_pcs[7],pcs_avmmreaddata_8g_tx_pcs[6],pcs_avmmreaddata_8g_tx_pcs[5],pcs_avmmreaddata_8g_tx_pcs[4],pcs_avmmreaddata_8g_tx_pcs[3],pcs_avmmreaddata_8g_tx_pcs[2],pcs_avmmreaddata_8g_tx_pcs[1],
pcs_avmmreaddata_8g_tx_pcs[0],pcs_avmmreaddata_pipe_gen1_2[7],pcs_avmmreaddata_pipe_gen1_2[6],pcs_avmmreaddata_pipe_gen1_2[5],pcs_avmmreaddata_pipe_gen1_2[4],pcs_avmmreaddata_pipe_gen1_2[3],pcs_avmmreaddata_pipe_gen1_2[2],pcs_avmmreaddata_pipe_gen1_2[1],pcs_avmmreaddata_pipe_gen1_2[0],
pcs_avmmreaddata_8g_rx_pcs[7],pcs_avmmreaddata_8g_rx_pcs[6],pcs_avmmreaddata_8g_rx_pcs[5],pcs_avmmreaddata_8g_rx_pcs[4],pcs_avmmreaddata_8g_rx_pcs[3],pcs_avmmreaddata_8g_rx_pcs[2],pcs_avmmreaddata_8g_rx_pcs[1],pcs_avmmreaddata_8g_rx_pcs[0],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,pma_avmmreaddata_pma_adapt[7],pma_avmmreaddata_pma_adapt[6],pma_avmmreaddata_pma_adapt[5],
pma_avmmreaddata_pma_adapt[4],pma_avmmreaddata_pma_adapt[3],pma_avmmreaddata_pma_adapt[2],pma_avmmreaddata_pma_adapt[1],pma_avmmreaddata_pma_adapt[0],pma_avmmreaddata_cdr_refclk_select[7],pma_avmmreaddata_cdr_refclk_select[6],pma_avmmreaddata_cdr_refclk_select[5],
pma_avmmreaddata_cdr_refclk_select[4],pma_avmmreaddata_cdr_refclk_select[3],pma_avmmreaddata_cdr_refclk_select[2],pma_avmmreaddata_cdr_refclk_select[1],pma_avmmreaddata_cdr_refclk_select[0],pma_avmmreaddata_cdr_pll[7],pma_avmmreaddata_cdr_pll[6],pma_avmmreaddata_cdr_pll[5],
pma_avmmreaddata_cdr_pll[4],pma_avmmreaddata_cdr_pll[3],pma_avmmreaddata_cdr_pll[2],pma_avmmreaddata_cdr_pll[1],pma_avmmreaddata_cdr_pll[0],pma_avmmreaddata_rx_dfe[7],pma_avmmreaddata_rx_dfe[6],pma_avmmreaddata_rx_dfe[5],pma_avmmreaddata_rx_dfe[4],pma_avmmreaddata_rx_dfe[3],
pma_avmmreaddata_rx_dfe[2],pma_avmmreaddata_rx_dfe[1],pma_avmmreaddata_rx_dfe[0],pma_avmmreaddata_rx_odi[7],pma_avmmreaddata_rx_odi[6],pma_avmmreaddata_rx_odi[5],pma_avmmreaddata_rx_odi[4],pma_avmmreaddata_rx_odi[3],pma_avmmreaddata_rx_odi[2],pma_avmmreaddata_rx_odi[1],pma_avmmreaddata_rx_odi[0],
pma_avmmreaddata_rx_sd[7],pma_avmmreaddata_rx_sd[6],pma_avmmreaddata_rx_sd[5],pma_avmmreaddata_rx_sd[4],pma_avmmreaddata_rx_sd[3],pma_avmmreaddata_rx_sd[2],pma_avmmreaddata_rx_sd[1],pma_avmmreaddata_rx_sd[0],pma_avmmreaddata_rx_buf[7],pma_avmmreaddata_rx_buf[6],pma_avmmreaddata_rx_buf[5],
pma_avmmreaddata_rx_buf[4],pma_avmmreaddata_rx_buf[3],pma_avmmreaddata_rx_buf[2],pma_avmmreaddata_rx_buf[1],pma_avmmreaddata_rx_buf[0],pma_avmmreaddata_rx_deser[7],pma_avmmreaddata_rx_deser[6],pma_avmmreaddata_rx_deser[5],pma_avmmreaddata_rx_deser[4],pma_avmmreaddata_rx_deser[3],
pma_avmmreaddata_rx_deser[2],pma_avmmreaddata_rx_deser[1],pma_avmmreaddata_rx_deser[0],pma_avmmreaddata_tx_buf[7],pma_avmmreaddata_tx_buf[6],pma_avmmreaddata_tx_buf[5],pma_avmmreaddata_tx_buf[4],pma_avmmreaddata_tx_buf[3],pma_avmmreaddata_tx_buf[2],pma_avmmreaddata_tx_buf[1],
pma_avmmreaddata_tx_buf[0],pma_avmmreaddata_tx_cgb[7],pma_avmmreaddata_tx_cgb[6],pma_avmmreaddata_tx_cgb[5],pma_avmmreaddata_tx_cgb[4],pma_avmmreaddata_tx_cgb[3],pma_avmmreaddata_tx_cgb[2],pma_avmmreaddata_tx_cgb[1],pma_avmmreaddata_tx_cgb[0],pma_avmmreaddata_tx_ser[7],pma_avmmreaddata_tx_ser[6],
pma_avmmreaddata_tx_ser[5],pma_avmmreaddata_tx_ser[4],pma_avmmreaddata_tx_ser[3],pma_avmmreaddata_tx_ser[2],pma_avmmreaddata_tx_ser[1],pma_avmmreaddata_tx_ser[0]}),
	.avmmbusy(\avmm_busy[0] ),
	.avmmreservedout(),
	.clkchnl(chnl_pll_avmm_clk[0]),
	.hipcaldone(),
	.pldcaldone(pld_cal_done[0]),
	.readchnl(chnl_pll_avmm_read[0]),
	.rstnchnl(chnl_pll_avmm_rstn[0]),
	.writechnl(chnl_pll_avmm_write[0]),
	.avmmreaddata(\avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_AVMMREADDATA_bus ),
	.regaddrchnl(\avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_REGADDRCHNL_bus ),
	.writedatachnl(\avmm_atom_insts[0].twentynm_hssi_avmm_if_inst_WRITEDATACHNL_bus ));
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .arbiter_ctrl = "uc";
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .cal_done = "cal_done_deassert";
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .cal_reserved = 5'b00000;
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .calibration_en = "enable";
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .calibration_type = "one_time";
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .hip_cal_en = "disable";
defparam \avmm_atom_insts[0].twentynm_hssi_avmm_if_inst .silicon_rev = "20nm5es";

twentynm_lcell_comb \avmm_waitrequest[0]~0 (
	.dataa(!\avmm_waitrequest_write_int[0]~q ),
	.datab(!avmm_read[0]),
	.datac(!\avmm_read_r[0]~q ),
	.datad(!\avmm_read_cycles_cnt[1]~q ),
	.datae(!\avmm_read_cycles_cnt[2]~q ),
	.dataf(!\avmm_read_cycles_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(avmm_waitrequest_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_waitrequest[0]~0 .extended_lut = "off";
defparam \avmm_waitrequest[0]~0 .lut_mask = 64'hFFFFFFFFFFF7FFFF;
defparam \avmm_waitrequest[0]~0 .shared_arith = "off";

dffeas \avmm_busy_r1[0] (
	.clk(reconfig_clk_0),
	.d(\avmm_busy[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_busy_r1[0]~q ),
	.prn(vcc));
defparam \avmm_busy_r1[0] .is_wysiwyg = "true";
defparam \avmm_busy_r1[0] .power_up = "low";

dffeas \avmm_busy_r2[0] (
	.clk(reconfig_clk_0),
	.d(\avmm_busy_r1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_busy_r2[0]~q ),
	.prn(vcc));
defparam \avmm_busy_r2[0] .is_wysiwyg = "true";
defparam \avmm_busy_r2[0] .power_up = "low";

twentynm_lcell_comb \avmm_waitrequest_write_int~0 (
	.dataa(!avmm_write[0]),
	.datab(!avmm_address[0]),
	.datac(!avmm_address[1]),
	.datad(!avmm_address[2]),
	.datae(!avmm_address[3]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_waitrequest_write_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_waitrequest_write_int~0 .extended_lut = "off";
defparam \avmm_waitrequest_write_int~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \avmm_waitrequest_write_int~0 .shared_arith = "off";

twentynm_lcell_comb \avmm_waitrequest_write_int~1 (
	.dataa(!avmm_address[5]),
	.datab(!avmm_address[6]),
	.datac(!avmm_address[7]),
	.datad(!avmm_address[8]),
	.datae(!avmm_writedata[0]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_waitrequest_write_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_waitrequest_write_int~1 .extended_lut = "off";
defparam \avmm_waitrequest_write_int~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \avmm_waitrequest_write_int~1 .shared_arith = "off";

twentynm_lcell_comb \avmm_waitrequest_write_int~2 (
	.dataa(!\avmm_waitrequest_write_int[0]~q ),
	.datab(!avmm_address[4]),
	.datac(!\avmm_busy_r1[0]~q ),
	.datad(!\avmm_busy_r2[0]~q ),
	.datae(!\avmm_waitrequest_write_int~0_combout ),
	.dataf(!\avmm_waitrequest_write_int~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_waitrequest_write_int~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_waitrequest_write_int~2 .extended_lut = "off";
defparam \avmm_waitrequest_write_int~2 .lut_mask = 64'hDF8FFFFFFFFFFFFF;
defparam \avmm_waitrequest_write_int~2 .shared_arith = "off";

dffeas \avmm_waitrequest_write_int[0] (
	.clk(reconfig_clk_0),
	.d(\avmm_waitrequest_write_int~2_combout ),
	.asdata(vcc),
	.clrn(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_waitrequest_write_int[0]~q ),
	.prn(vcc));
defparam \avmm_waitrequest_write_int[0] .is_wysiwyg = "true";
defparam \avmm_waitrequest_write_int[0] .power_up = "low";

dffeas \avmm_read_r[0] (
	.clk(reconfig_clk_0),
	.d(avmm_read[0]),
	.asdata(vcc),
	.clrn(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_read_r[0]~q ),
	.prn(vcc));
defparam \avmm_read_r[0] .is_wysiwyg = "true";
defparam \avmm_read_r[0] .power_up = "low";

twentynm_lcell_comb \avmm_read_cycles_cnt~2 (
	.dataa(!avmm_read[0]),
	.datab(!\avmm_read_cycles_cnt[1]~q ),
	.datac(!\avmm_read_cycles_cnt[2]~q ),
	.datad(!\avmm_read_cycles_cnt[0]~q ),
	.datae(!\avmm_busy_r1[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_read_cycles_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_read_cycles_cnt~2 .extended_lut = "off";
defparam \avmm_read_cycles_cnt~2 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \avmm_read_cycles_cnt~2 .shared_arith = "off";

dffeas \avmm_read_cycles_cnt[0] (
	.clk(reconfig_clk_0),
	.d(\avmm_read_cycles_cnt~2_combout ),
	.asdata(vcc),
	.clrn(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_read_cycles_cnt[0]~q ),
	.prn(vcc));
defparam \avmm_read_cycles_cnt[0] .is_wysiwyg = "true";
defparam \avmm_read_cycles_cnt[0] .power_up = "low";

twentynm_lcell_comb \avmm_read_cycles_cnt~1 (
	.dataa(!\avmm_read_cycles_cnt[1]~q ),
	.datab(!\avmm_read_cycles_cnt[2]~q ),
	.datac(!\avmm_read_cycles_cnt[0]~q ),
	.datad(!\avmm_busy_r1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_read_cycles_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_read_cycles_cnt~1 .extended_lut = "off";
defparam \avmm_read_cycles_cnt~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \avmm_read_cycles_cnt~1 .shared_arith = "off";

dffeas \avmm_read_cycles_cnt[2] (
	.clk(reconfig_clk_0),
	.d(\avmm_read_cycles_cnt~1_combout ),
	.asdata(vcc),
	.clrn(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_read_cycles_cnt[2]~q ),
	.prn(vcc));
defparam \avmm_read_cycles_cnt[2] .is_wysiwyg = "true";
defparam \avmm_read_cycles_cnt[2] .power_up = "low";

twentynm_lcell_comb \avmm_read_cycles_cnt~0 (
	.dataa(gnd),
	.datab(!\avmm_read_cycles_cnt[1]~q ),
	.datac(!\avmm_read_cycles_cnt[2]~q ),
	.datad(!\avmm_read_cycles_cnt[0]~q ),
	.datae(!\avmm_busy_r1[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avmm_read_cycles_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avmm_read_cycles_cnt~0 .extended_lut = "off";
defparam \avmm_read_cycles_cnt~0 .lut_mask = 64'hF3FCFFFFF3FCFFFF;
defparam \avmm_read_cycles_cnt~0 .shared_arith = "off";

dffeas \avmm_read_cycles_cnt[1] (
	.clk(reconfig_clk_0),
	.d(\avmm_read_cycles_cnt~0_combout ),
	.asdata(vcc),
	.clrn(\avmm_atom_insts[0].avmm_reset_sync_inst|resync_chains[0].sync_r[1]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avmm_read_cycles_cnt[1]~q ),
	.prn(vcc));
defparam \avmm_read_cycles_cnt[1] .is_wysiwyg = "true";
defparam \avmm_read_cycles_cnt[1] .power_up = "low";

endmodule

module wr_arria10_e3p1_det_phy_alt_xcvr_resync (
	resync_chains0sync_r_1,
	clk,
	reconfig_reset_0)/* synthesis synthesis_greybox=1 */;
output 	resync_chains0sync_r_1;
input 	clk;
input 	reconfig_reset_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \resync_chains[0].sync_r[0]~q ;


dffeas \resync_chains[0].sync_r[1] (
	.clk(clk),
	.d(\resync_chains[0].sync_r[0]~q ),
	.asdata(vcc),
	.clrn(!reconfig_reset_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resync_chains0sync_r_1),
	.prn(vcc));
defparam \resync_chains[0].sync_r[1] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[1] .power_up = "low";

dffeas \resync_chains[0].sync_r[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reconfig_reset_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_chains[0].sync_r[0]~q ),
	.prn(vcc));
defparam \resync_chains[0].sync_r[0] .is_wysiwyg = "true";
defparam \resync_chains[0].sync_r[0] .power_up = "low";

endmodule
