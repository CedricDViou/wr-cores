// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c8RhuH9YMzgh4Qxm1hmVUSTq8Blq7Nx9YnmxS0rJX0Xu/Waw4UE6LUi/VgPkAMsy
vmxirDPb0HKNNrPOy+uEb9fItQLmUyyHIBo5CJo6MwbLkfnp4W/0em9W7N6GIO8Z
pOBUjtg/g0R8vUQWKrR2m/OCzUJg1rR+HE8iUWeLuos=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6224)
Ktk28l0rI0VoFiQ7TiDc9ZRQiPdQ9gNs6/EqoNq3p/gsvEDQPEYxLaYOY8EMJJde
/RIrdGOSuufsMrMwcytXVQs2yjRMfeEn3Cry1KBbPW5P9vXMZxqYL6RC6EA0FPl1
ig+Lw6Q3/hPWvT97u5iyEPzXu1YGz2oS4HcSW7wpMBne6c/XM6Ivx8TC9dhY7IlT
9PlHKAGrdXneF+MsgHKuMjqgYPSNkiRELE5ywX8SgFN+c+D/2O/L+DUi/zdv6Tuu
QpNepRma6XuYoY4Y6IFAxigOh/cNHub9Ujw1ozymTjjGCNzNUQIbHM8C5ebUg5OZ
PcYh3TM+H60T8dQTiX+pedSwpMRSj/FyaYNpGReGQD6pEr10XGesQgcO1/viR2Fe
9KzT7iYCcKdMZ6uLa8y90VLIl3ycaL2W/bQA/RlTTudBJuAXi6WlH6Yl7a5n07m6
k0JZDHmt/HzyWDy9vYSWuZBhGpN8Ym59OmGiiMuPTqp8tUj3O0eNAj1J+KUEXPqx
wJW3dYQorZRmxDnIljS05n6T2U1beKtj+HMr2zAj1r5mNScHqOMgGKi5zENY7EIV
+2hv4tOxpYIq/Xf1Ph+wjYUDUncFk9seX19bkSg7dCiaJPioIXAZV0pnYc3++Cua
7slnCHPOk3pda6s5PCphrSdbOj4RH6Wv+LdBryxUssBxA6R55osnwbSNIX3Brw+n
iIcHqswsPJ+Ca12+mBUEnbaacPqFcjenEOSzns9rVxKyLoZaycEcR74wH6lgUlRN
OtglZ9NFiCBxlYgwB+1oMaQ/MM+GUWQtbcRv9QKK6WaWi1stzezryrdNbXqtsUT5
+MjlQNkcJou4F8haw4I+tkEUIydQyinPykEntNtt3CRerOFrBIu0qBgyehQEgrSO
jJWm7bgtGMUSKs4nxXTarRDf6XR+mNChE/2buKqO3TOLLB/EYefvEqqxpBa5owmo
ylnyeu2/pDPlHc8fLma0TnwMFbiuaPAK1Ngm7u0/oBOW5mrQdh4kN4LA70K2tNlv
LgjlUZjSoXuPYhDafT4tvxvgn553JxVfwda+cdydo25OyRGStXOkbz/Vcut/pbQi
A1FEy3ICECpkKPAkLEGu4wX2ukygBPyosVSxL/rD9oggSaziYGT9Na8i0251zzr3
y8S9XDxRVOPlyUc3E5QbfIchthjHha0+CmfMRGLPu12UGu+DLeyTzKS5p1HeKYiy
jdy21LDciOuhuY19+doSpBHGqyf0d6963Xc80Yv2+Sgxov8WPt388q+bk/a1di0+
Bz4z70VrluyuWovnAvye7ZDIZcJjzCvuszqHe1lv4KRG9Qgz/WTxtc3vKWwHnnZ2
6DIDADgoR3982NijgAge+l0XuC3TjJMdH0mMHMbrU0nI6nT7eSzsdgDnqAL5KGFy
nSi4lPuKqlGIblxW4S7izTHaES1SAk9sN3MQLZNySimzkgU3M8Cfwdp0pUuEyCOe
3hYMbem2mKiwkE0P1PNn6hvq0uLRIQSyW34g08bIB908bLUBcAyLmYNiv2W+wkIV
RgeSsmq+XrsXIoxwmhfCWXmh7Z3Dsyo4i8XaI+6VODxeXU6kE/hX+j9X4elVYvKp
9iKllPuUjFNLjShsQN1QDJp2E4MYBv8gth83x6/dH/t57G10r4/G9oMsKyzQAb1+
aViZeKJCLhFwJB9L4/3FL4cZMaZMe3qMiUs6ydRTNRBIhUtZNs+vUaeD3cA7Et3l
jG+2yIgyQ9Zm+/7XwDzPLnrkOgjx6Tf1HQSeDN87Ta/j9ghp69/Y4OyN+33HqFLx
FXvhlWd5FmHeQ9dySf6feaKHwg9yLLgueysoCkfM9kxd/AFSEc2vGy2fHZUrlRi0
vLtlTyJoumeHwmPesF7pgF6J2XWTCM8UnWvNv8GSjvONFtMJrMTSoCW/lV6wXaEL
b3UyAnjViFCoyPIbaK8L6bY0xXdMpScrgIYPj26fQPjitiiA7lsLaagp5RZF6WSl
WaT8lRTjGk+hOIS2ukd/QBsRqndmh5t5EAlqjhriHz6FSmJwU3vg/OKfha0W1SEw
pZbvZ1YqtNY36/96J5o30YWElcYMAm9Z3PlhoM/h3PebU/rf3PA5vGw94xtcvmt5
Hy7WMIE2pr7VEXbPVBmuqtumuISjvFFOhLvfInayN6YJ/sL7qZQzahOKK2xwX5DB
KlPSUt3Dizkp6vwp18V018fpNfEeBMwnjMKti8jZj5fS1VpXG4VWtscQrc4Vc2IE
pIN849uvD37jHjad2T4kvpGbSYO4O5FmxyQmLXXu26roA45NRsPD3D+n1ebBKpQM
8yluDV23V3q0qjzy4CoBwswZEwiJmsg0tUilM+ha1/ak1L5d4mhw8pxzGX0ioj2W
mujs15CjwpiiSyXY1JjSktSOE/eeguq/2C9Yj8mRkaeTJsL4CuTUAFNxw94gAx0k
I/3TIaHn3Juk/jh7Zv58Mi64yPGkYg5HwFABQcAU7I8mzPSbuZHvsiEPfYw7yQYr
Q2y6tvRNRMBDJN4yjuGpHrHLhf4jZIttPuJu+TubaGrFGZMloTqzlY1GjJZ1aQJ0
vYFxtkgPsJYw9ttgdp+Nd4+pPdyTZNkfM4IMN7Mkkv2Cv/UjX/ZUTjMr+erdjYJ8
RilkBDumbcxoPaVLo53nWTlFxVTOynAHrHIbC2AbzOzhnUYxFLXq3uqHk7VevnwY
cDT1pJPcMH7XxLZy5tfII9PXNbACQDkZob9TpMeE4mciXXWP5lQypKn5E6gdy04/
lbYbnuylOB6f54E0DSJWhPdE0Xrru49eBBrQSiWjjnu7VqlE42/1X/acEsDq3iSA
X6yE99zA3HIcsKyqvcrk62kf7ZkJgSO9cdIy3AXie66Ul93qOrK3Wc+2XLpLniO4
ESBLlTTWYwOpFZOLWfXFXxsSh6ngBSr8hlibAOzV7MJ/8YFXvHQ58+lTDEf6l4NU
uVFS8zBlRXFHrMre1GNZtgg7969aQYv5SVl9fph1pISQ0Y+F+HCEmU9Oy79HL4t2
phmd5T1XPQ2k7+jTpX4ymHm0/JxA8ZrIJxBzknoCVyTrLC8F/p8p0N2A/Hp0PLd1
waVw+RsJafZZn7JO5pIAZ1cx+1Ul+qUHMzt28PZ9OlDDBuZGFAFaASIx1T5xMS1a
9CKmUvjrUMCDnsDPYYhYVbfcfIwnJvCAbb2yMYGkTKYcIw19t61cyo7u1590kmAZ
C+TDPXtSKgg1vq8A6KAnZPDoz9mXPRSU2/q9WP4kg18bowabQlpHeGpGtqRK/AVp
5w95Kf6eFBdt6mxLk1DZRm+51d7VsA+nylMnY72igvwpFaqREvgklOEQu62mt09+
Yu8Kop7HEMdyBZYZv58CjajyOnHsBYcBeO+EmZnaTfkEeQ+P8RB8dLc6WsVy/vGw
RBzbGHFNabWQpqFxHO3cxBBpE3Flb7moHbiCB8avnq+9p+fJUmB+n1rK1AE7kUx1
tsegAWI6la8GTpt/L9arsNOwZ3AvBs0RQN1RwWuS97ujmJ+5qn1Fs8Mw1Bweg4RZ
zO3ifetLAQMgDsj0X6tDCwe1MuyIlG+pcrIdFA3O80sFFM2kCuwGahLLLNm+p3Ff
+2ceSr5FFBaxbWib6rHhacPrkMXxp3yma+O2BRc97008IaFzE6rhLcT+BFFfbh3V
aWxyIixq9rWtJYHVbQwKPy2u0GnlbG705rR9815DILI358eKmP+xyRqHOtOgm2Aa
mRaAV1SXYZB+MW3A2QF4hO0aztt1jnxNn2TRDreEP7dJ2CEDVA4cn9SV+AGPGFwM
0EUjwyrclFxEV/sF/cQjc50onCOkne6wYxpe6wJXi0f+aT6a004N5r1EDMX3fCI3
OXIZnxtsTbDM+2LnNUnM+e8bLAV5NVyss2ce3vslKXkhPYBxKqVAzk9vMdCVG+CE
RtOTiKfQtRWt7uW4q46lq6PxDNyDcFuyvm58SK7W9hCxDGkiQivSivxTaZ4u7IiT
+2Pk/RIQb/o9hnTjXx3sw+c95Ewzrq3gIdSZSukzyPx9RWFOC3nu808RO/HbHZsG
lKrhtVJ/D91lYPc5CC5OBwqhtLd1yCbqae4aZz0BKcAPLQ1ScPVxY3niDGs4FdhX
spJzxL0eJEF29nOkke921qLzb2oUKIQJ3gWL6iM9/w4UeaBc6tLBIJ7W8t76eQj9
2ce1dirjTMJdta4JCaToqoQV/dMOdBLGnZ/fougOKVRpmFzAJT76+PdbcDcDYrQV
gBfJzbpTadMqfErvKoGorue8eBUm3lI6Jh/LtB3QnPimkWLDuNWXf9GlXkNeVsW9
48x4m++NuipUWW9J5/UeOx8hogEy9z+hGrw7biDEjBPw5qh9VvAcmz6l3hdAqcQW
YUEzAUul9PfPfaj2whwTJL40BvTWC5cUVoJ/yn5ev4c7k/23l4ZBAkzVFbQtYs5c
k60Oc5sIqbVLa6aXOENfpB5Ba3ADZR/SKaEiUJ4WBj2iob9RoofEF4mKaBTQG6GJ
A3oj5uqUdhp8tvZv2VQ6Y3hjqrnK0dR76swmsc/K6zBAj1CWmMsEztnL0JJVKGFv
u7wFwqsr1UP13UoPrgCvI/ZIm2GabGxMKVLG87jOprcShpiNX1t+Zn5jFyy+xBtg
kUcDrKA6NTvn+36BK2LsKBxLm8889U98IydV1Jv5w14xyEpFilm2A5+yWazsw8mO
VOO7DnjRlylH6Lirc3p0uzQNFNAFYcJ3vq8OyW2kUvFN2JXFde9fGHRHY2ERxP0M
rqNiqluQIa0AigTCLjFbk3R50hQkCkfXyTbBRFDQJscmRaB2yLco6JySvu6+wdsp
5z/nx4MvaQAFxlNm6C6s382KXylno4w92lqNE3P6KgRijgCBMFzygqSdtjeYY15v
mU7e9S6pInH+N9bdawsXdJQzKABv7Bw2fLOkZHBCBfIxNTasPA+QWzuvTZoS0MPv
QhXBoyHLt41thWQ/nPSdpc8GHN8nqg2sDzLSif1hgg7r+JsVMCn5LrCNVG8AAX6m
Syql9vHpSRCPBD9CYKgJ86beGTxcUfNX6E++iizv4eKyiJ5tXgLZMSL3fA29Ybcv
gjVHwAa6K/IAT0su7vDeSgBiS/vaqu6YVYl2BYLectwSzIDmBabnOjPxhnfITTdb
2xHRKFxPT+fzSrPpSAhrWHoTbw4t0QqaTELtOuY8+PtlKXWAXryr2UYnauvDFBvE
BZ5zmoc2BVA4/WFBD+CJNhuv9o9qN03ZlQS5weX+aUym2TtE6Tw5MTToheAN7CDv
r9Co1wf/W8cmFPaiV3xzoDDaw8/qMlO+GWCg18Nv90v78zZvKaj+7J2DDDcNB1iw
XUakA0yqdE2DVaEWDTKXtc15Ybz70tJXJtu5kyBkwKCEG8x6h7QmKXVUTi3adnVP
0xrLoeQ0R4DlOvwa3f6IATOXEMKdi5GIdf7guaD7PlpUbxfAtMbfUquwxMQu2xl4
47KYK34x1X3s4iZGU6iC5evM4oWlM1JKVoQghDR7dalfoqDzzUhwc73ZLOHPFl1D
aWw0wrMCAHTeUVXwFvEiEkPBbUtCVOn5tOYwkJ0dbqdxn2KpNXgT/BZLejzyL4nO
xRM88va9Vu1CJPCz3a7FQWPw9qdBAcOJEcOrZt3QhrzI+K2GRyyB02XF+CI6jLaK
Bgf465Svm3LLI7joEU6jkp6V8svULACGj+BAUmwAkU+Tv+Of/3Tc2gn5SIiGPF69
5Rjvoj3oWzO4XVyD/8LuQgubS8qZbn4hxDzgb6T0w1NhM7XJMJzUDwwvywCuEYDc
Q1TLN7jLosIxwKu4Blx3HJPxpVYlfs57hupZhPN20IYl808peIAwdI/gRJXB1rFm
zkr/QyZXWIdf3eg5Mej7LBmymMkHWLGjF5GoiHzpH6KF28m3F490Uikdfcriyo/B
IZBVjx4wy/DSLmLWav/HNXyMEeeFxCoRPkAEykr2yh8SdEhKlACxibGq6xT+mSDk
QU2N/f/J3G2M4pB0paCmQXbARCxrXNouDjuppGMJaWYaVnJpBe1auOLWpJdhmdSE
RPJoHbzuDgw+6yY2HdvF0dcmuyEt0hU4xiSbVopd0sSV9sffkYr5iOZg9rDYVRvi
LmdA/FSAOLg4KyaO1T47xdBWYJnYngVYucH/1YC+J7UFvzDLNsGnq4uqa3xIVjqf
Y2eO9sbzjzc5FSSac4kJaGc5EscxaoYqB1B3SMAm6AkEjkhrj/s3Lxxfot4q7gDD
ojWGrEH/+Ba3knppNA8nmTUlYgR2fNuWg6kqmuJyz92zVhD8TSKXn3OtpPqxATle
gcuViqwaPJuORkS7Jq7y8Nu5pgnnF3ZzKOUxAR9KnODlST1e3BgGEtHiTp/9StuE
VgsN2JNOH5+puqkjI9ikaKm9p1U0DnLghqY+qEe4fbq+KcpvjI7bsrlyj5oyr5LZ
FsgXIwiA23uTszsDLSG+kRft90tOGu2ZEq3CdXu6OJ82XP0Ijon+vhCHVjWcZHor
R+T3iy1SfYzrAcRIQ1jae2AIBsU9xj5i7tecvXDL2haBbTOspkjfheGT94JC/XXf
MAHHROkZjWFFflumZpotlimDwEkDa/p0yFbTOg52GhNK2sGyujt3/ke8wnQj6GKN
3qc5vTcJb/RZivimUl7EOh1MNHDZtE/TEdJTDomMqHcADbgwgnUyYwzC0/2rhGl6
YZ4SmsZI92VJp6/JT0pTmKSHzTVl8j6kDUtrclWpCSW5G27aNhKcm1z5EH1BtsYd
ZslbBBo1yleM0ZKhq/arC27EeGYFnlIjWloXuSveP1P+dh+9u59ucuuoBMCe1BKd
1kO1gKEmu88R/QE86mKSc73NWaDAIPQ708t/jPayLnfQCIXolAMUlYT6JqG08fAk
757CKKenyrk9N5tSE3uI+J6e2zbKBCkL+sJxMjQnjQ/D38KdlgdOABWgniHHjFAE
0/Db6DolvtrQJUv/N8S+QyMqhfNXokCsLSjRybwDnuqnk95sMmSlSaYAy6cToYvA
3gMYdmhkJIWhTvS9yelrg9LiCWoCq6vg+MbKt/P7iVtAd5zgIYBQFaAlshZH+RTB
325tv+rn6f2vludwLiHgwlqXStsXZb4SO3E1uCtC2e16sC+b29vIMOSaKzwkVgus
FMXxK7j0czCCA7lfVqttTNLdWLIW17Zn3z7c62ktqVJZOQIcWWOz6XeBggQwOX3g
/JC0UpzyhAjvLxS6fswc+WC8iSrXT2mGF3q6Mox5236CWKSuW5q/QkzfIk3fuH0z
Oltxppf8tWU6OyEns6WUyYCY88UlbyQ7l3TDH5qrCSGiFcZc/6L1/TkNjUfvtTTj
o2mlCHTHVTbHa55qZdCdjMmN3oK1yfNQBJRqkfVl2SS628lsSMb3PryTViCNMkkM
zLJOd4s5Zrv3u1IK2zZuiPA8MDOfjZ0C/gUhdmoHIfaleu2qL/i2SK/RRoVuRgfF
MWHIhx2fbVLrmA4Zs6lRZZjkO+qvtZTxvV8onk8aI13N3L4CMQ8W/AfnvU4wn3yN
jkjH3xqMOogNF5uwRH49KNUAljWxPc6Qe+K9dz7aJ2kyrtVqXrxeo0N7BNz+U3Uw
x8eaF3cJwiuEaK/TO8z3rtipR5ENBm2JYwo580N7VfpaFki/2xdjejWRVfKPb02e
0P1l/GaN9Pk0Ar/gdD1sZofik23zuF8sO/UOgZNEQ376nMSJzzztFY8qrRt4cD5P
LZJGd37dJucnZp9BXccpRYTCFkrwOdalnZZtCEUtlQyPkMgY4c8fFBbSHoxsMZe0
34rXueVp0UPfeCKf9FsaTkAMWF7TQ0jv7QiVh0i1PfKkvRNAFmsah8SKoqggjo0t
l/fMAonagUqOl4E1uToZ9vwUwVoq4Y+zEkpn9PkH1DGzPk/a9BCeEa7puyOy33fk
/M9V4MW/mBJirlPe1ssOySG4oLoZmnjmtZ7nSgPzZ/pPpKVQrK1X1rOUjZ0Xo/US
NEDSJozJdwjfJjpqCDKQ1odOMNxb24DoonliYRoy2R+58nih3QXEq0gjB3ThnlYN
Fszx9ZC/HRKh2cd0raxpiXFwDn/M+qgcHYXQvADQxrKlPNwVI+LIgWu6AH3o/upG
o/1VDi5aPyZThh0LUXAZTgoaBC4g6n1iSYBMuuQhgZmftTSC5J2e1LcjsTWHUIRb
tCegW8h9Y1wC20YGFzIDF8gIvTg+QtJE4MrorLG9vBsIJpCDvQ3p9v9uzt2TGNzO
mSf3Pg+Ps4Omvj/E+akRNO/xuZPJerdJ/b0jYPoOFb8XCR7U+qrecS+WFb6BdtQb
jnYaDUOxAwP9S3abwXBP6mErw676azwDAhGX61iVkJw=
`pragma protect end_protected
