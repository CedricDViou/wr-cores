// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
agoGW3xt4dSVpsyHkNHnkCeLyT5ClR+O53KTWeicCZz+jfJ7oVUbOegrXUAaHkKJ
B9YFUQLtU2E46yDLmUcbZliQQGZsd3D2+cq2jojlBlrE8PbFRzgGP2242HRYyuIO
VVS72KNWbtESOMRY72adWXYBPLBYnekJaC5L2dGq9U8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36352)
/m7IuICmevryWBvGVjQEl1fP+D7n5kfDcSXVScAckdqi+567ykMyMSS6m6dMUBPq
bTo2lump09DWbu4stVwmuRD8/5l4oiy398Ooja2XJgw9rx8NS/mBTU7O3fprub7S
y1WNtiQGsepzF0Q0NgK0JjDH7KISbN2DlV45zGY7MshX7W1TcI5717X2hCLZexN2
/iGkKLDQkvIJSwdjY8W5IjRHaBK1FTaaqxFD6j/eOHeO16VhvF9fSVcfmzRBkhhV
jIIZCNl5nHIkRYCR9qlhRuZYiGwSvjsCZPWrgsnY2huo4oHDizzk/GfHEqBTSEp+
74hh5l4hH0fPYn2b2t+mktAQe1Tr7KXfPpmw6EIpmm67ZqHprfyxhn+bn8lm6ADJ
sdo5GCFakXtBq/Vq39VekYuUb/Q/4ecRd5cQutjgf7FfGrLY8IDNtOvr7rl9QGUj
wW5eWFWSRdBKiTUPMjEN7ePl3mTL/57/qzn9qPltNZ3SAmFudbShHuOtjUkz4aFL
CBt42bsLvDyjfLc+ZRRHqA6S23i+ABTTLKU3glvnPRu5fFGGsny5xn/zssoW2dbi
BZIPDZ3SYwiduv5BSMWrUGC7EqyDk2phL57sbZJDqWLnjujZY2y0DxuJ1G+fSfdA
VjEDeybXc09Q7U5ASXNlDNs5yBYsu9f9G673EFpXkG/0IHX2F/sfu4x/QZC7Z4bX
PpPlGO+DOPaeB/TycuUdkfXK2gHM87Hzl9E+suP0f8/tcePmeZ0jLaeLuAFsntS4
YvG+nX6AdpNhbXV4yoAOA/Z5mh2u0pRiom4QSlNKpNmsZFg4PrNS+j9M9urFZ4hC
c00lpO0twmto3aoCgCMew3wHsqywLYdvnhtTvwQLQrr322ZMmQZywYIM/jexYwR+
hNkO92HWZUOsiYzFvUdm4jfw2pFjYOLrfVKBL4vPpohg8WL6znkKt5AaDOQKG2gr
VIx+AaqZLX4D5HrWZOjszuNMgmcmITbd9pdoejnBxFjinPFrIjAywx3nIk59dIsZ
SMSzFZCXsjK2CViplDcvbpqxB8MbR9eJ/csJfCpMwB6MGC/HpV+bxvkg17dbjW1P
SmdioaXKUce9UC2srcciviewZjivYrutFhhxoT2rf4gySASkSm3+OQsEKQOtpLsd
TBE47tb+la8uHTaJfPvVXC+yrqyBjIdfVn3HkjmWFjVi2r2rSvqEITbSLdpdDSfH
DlW1M5quiFQsVSjQUVF5jMoYihtd4sj88Fn5AjcARjNo3bvSuMT9zhoqRBCYK8Mr
u3V0D3IiazCKRPH2wt8ArQlUU8pWQlb0/sxhtERdB8nE7RcV0e8pwEYLUfuf4xT0
/1+74c+8BZRGFT+E5lGKDTmoBG2CHqwLWNzUZjl47Epofa81iptCmQPRdNRwT0S+
7ejhECUiCW6FPEy35qJ1KGfylwfX55xGsSoDOcvsfSGFQY59gSu7qF5rHX3C71NO
oVIzIw71WKINBtDlD5OQcUYEA7mjViAKEwemFDosmOen5XJpKDi0ZRTEXB58YqQQ
SQJFD8D9+2K9AIXxrT4oR5RPUyLT8EIxdj6Kz95Ehu82O8zraM6EBptV5l7Mx8oh
0JUsl5JO4SfBG3q+owpM3mF6+lAF8RDgoCk6yawE+af17zAMEiI60DajW8OK3RZI
1rpFYRRe7IXmtgq5lcL7Ma7Uosgu1+t8XRko4ZQzKRB0KGeDrHp9FygyBugm1tw/
yNo8RD++ZwcaU9uHW0pDzfm4o0+WVGqrEIPqEFLCS29Dnjk4gFwlaCSWi20sCPtP
S3ize9P78YvJ6e36VCyIUaNFL8W05oDPqnnWUuPXA+pfQTh7TJ3hLPbdSTg9Y4+R
3/irNYb1QfcAYTZWxRaGNX1J3j11UheYvNcYa6v7dr+b5CasDK5rY9ZGuEIOgq2O
rAufngjARUrhM4WELuo4By4lRCpr6OMABCiJ6BPIReaeFSuC0suwaGgGdN3hdvRb
3Utqnqjios19+8sORHvhSXiz40uVV06kCvPUoFtUfJhME1ftDiPcaAcJjr8fhpAA
LIdzUUq0hvDsGxSEkmSYHRoSt0q+Vl9xgebEpUXIHNraBp5rZSIbFFnvIwZk2Le+
rgESVnnR2Bn9KgvSK34Gq9sbS7p+ystiPlqihDgXwQXoQlhj+2HMFyEper8JkKF7
oy5sh7sy3ZIe2t4bC5jmI5tE0QI5LVZdBKcvPHX3lxh1brsENmYLqgtlPINPKLi6
aBa2iqXFM2EQKFk6yv1YMYOo51kSDlGdmqHoQ0M0/fLIltBuNJJ39VCEEwXBiPv/
bi3V5+T07jtXFW1ttRVpUy1K2sTeUlvkLA4oL0UzgvyDPpyMfGWpWJ1rWspdgG8k
alEcY1JUkuaW3rdyW0mqK1mozdIsvuEOj3Wk5yu9463zmQehDAZmWh9VixdKZehl
ZYlpQBSm7fb21ndg9czzo1lwXDa59i9dsut8skJBkbcQr1Djf25NtQPZ2IpSh5Uk
2dy80Pp8uEROuPW1DtJwcgRlrLA8bHltq42Wr54ZNDxXOEYiqaP3GM9V9/4zfbdc
Z7xXKmcQ9mQIcWHleLLladFARTOGA3499Ct3o6l6KbnHwu9PkZUSsMAQJ8qlMcpY
oFYhaYX2/IZA/dBhn/cDSfhl+0w4EECGbBXvVuqxUU3Z2hHaj3mg139MhUDC2Kcg
elnQ+g5GB+lFYF65AmQSn2k3H7z/7Ben2Ka2pNcn7MVzCE8eblzKmIzp6Qp3/EKa
W62sIvJcOJBwlPPsoVY5VP/BZ7tmXJpB7UVdeym+UXYFLPYupri+QaDYisXEMCy6
ZdyA7JfFWtB16F7fJPro+N+v9ftKpzUHs2M7Lw95UhXI+63ghCe3n3KiW9r0NRsB
1/2YBIxHQ/GNCPRZkB/8AQath1zYevcE/7ejUu5/Cx4VK+3nLQ/lkUg3/c837l7o
jC1hpz5oN+skmW1BIEJpOEdsiqKTotwShUgU/pw5GopGNWaklY9cbIydupACfsOj
igkMPhmw6HzNGzlnh4TWP0G8x55OqUCWDHZG9TgC1RwBcNDB4YIJMbNO2iQ+qVIT
H/2ClOaEJNwPJv7p5GRN7kuE3qPgg9mAyOl9Xk5isCcQXCNTyZSfWE3iAzHAcUr7
aO29rNBnk95IQ99B7vFPbmGiWECETeFko1gIWBcAb4ESUTd71R99JGQXjlWTk2f7
TcSgN9ATseoov6P9k0LW+2FSurGHdVgn2F/gs6Bu52Otw/InTmzNRfu622UBcg8Z
lgRaQOPaJISiDFyyh9rARCckwFHZsQ3LlLChhUrU3NsJY8dqUgjQKqdcCHEAHYEm
Sm9gPlpDRK8og5Xae+sOuvh843Co2ZxL/l6T9wTvVQgrO1Awqrgo9QKuHk2hgFkK
k4rS5rOSUNkrjPtP6EAMotKu2mabgcIW5O0XttOFT1rycsZdDMKgBPsRipqk9n/y
fCUK3cdSrxNxf3kVYni0n/4+NMxVr8onpgq6PnvbW0t0m7HO1Cp7X/eF6d4NSdva
lhWQuvbtaBmMnmnfmAxVa0JwiOCErK3wWgCOpOkO7cwimucmJ1CJPGZk31zxe3UT
XqFwdPKXzHVA1L4yv6YqsVmpDUWRC3oIslE0jEkLopyhejOtQLneEacL5TnhUq5s
EPR/zq13KF8glPH14Ip6YK/44evfkUqufJxfeyMeaf3g8itd69j5MwT3L9PqiJfD
qmNgoZwlErDKuvFNhtA/MH/AxM74yhVfRK9aZt0liND1GG1XFsDGxZhF5anwxXjf
vFUjFjGa/hyhZRiI9Ax76MCZ0FwCH9ReysoUV9GKvJfTcSfA8LPojCA1wdmZce/J
3EPdWIlLu95s96yGjBx/S0e46SkgP2MKTnUS1x2YBZXZQgo0QQomto4ES1nZqv/3
aDxIzWVbvap+gEbyYqfanHgjfLgVyQMp82WVY89Uu+4CsJM8cm28GR3sP5y9yULr
u+Oxw5dVbUQeCuLxHTui7qL287jlCtgeQzqambDs1MCYabvhMUdQrt1/0ESyWI9g
rxnM+ekYdeMT9+XggwJ7afcj4tw0d8/vWfx2HbiPpKT/QzlO0NDKSkIbmqlfzBuI
7QWwfwIHmOGQ681uXnzcEd0YBiPuthzw3hebtZWMjQDjlq4WsvKrgx43Z0ZzWHQ1
5xo+qUIlOolguNSQ8sXbK2eGTDp8qp1a0Ui/PVp/liFI1Od54VgEexFjErsx+AAL
e/G2XzayTdhErtCB/6L7tdY6S2mhRAauFJmY0EUgRU3g0itgYYPO7tlfT5JgYwo1
S0R/fn6OjMslxgx30zKODtBL7/JvkR95ic8xrtCs1IcsKIwhtKugY8WjTQSmJ+jR
c/7l2TuQQ/Ed5d9gcFY4WfAyoo+qfUwY02cAO6Jc+WApD8m6DiK09sn2W6pW7y6J
mKMp4lCYIVCrOzK6q06flkY0Vq3RvR3sEnlT3VrCgqNuPoa+0GrEPjcJQc3zzRJe
kgaCfbxdvItZIH6PvOWY2F/Jn2eNkFahJLfs+X0n1gTJ6iTDdfn8OseyU/WAN88p
7LQV0DithZ2bqk23+D5uwWvZmodonlsvnV7QU+T/N6qjV3dlR7KPD4r3uuV9aeDG
IS08hzmgv81/VIjhPcZG3TIYLR8L5vIBB/NXEt1CgwluFPFvtOgjmCurSRzlsUni
Aqe+QyBnbTyPV7fuku3jlfa8qu9LET6meA3XLnAxyjIjJchmN+Np1A2thZMDF51D
eVYdJxGtZM2F5oneEqX55XRU16B5Fr1NUizs/VCopMhzYhK1CBuNyvcNbGr36JIc
NOqMSGBDR1QwhI/DNFZS3ny2VOV0jYzD1ouICKMx2cKcs5GBR4pIc5rHEn/Qgs3e
KyfKpV1xAuDa6eZGg/Q14i498hc7I7Jzmg77EsQ0UYE+V+x2eGDSugrBGnhV3Pfb
QwQViMRmeKtq3Sf+wQpCapnNl/URsKVqG4v1/5b1jO3TpP2xBY9lemTW1N0me/C5
ZzXdxkIIxiT83u7yvkBDhp1EuqxcvqvWG8IfpTeaEhNOgqNhiJaERXv2BR32lrFB
w/+MyT2lS4ubkdiKxnaQBlfXwyTFgy5T0QmTNmGO57RWRE7tGwEEOh32pBe2krH9
q0r1zBIqKm6fibT/dJmI5sNy45Cq/A92V0IhEMH9uXHYx0Ue5PblRy0ZxmuzGQIC
vlYywe/juNWPGD3Fu6vHg3TIbGBtDlZVp0K34+MaqtRnflD3NRbeVWrzUxUk2zTp
+Ddz5fVsjq1ySPE+arWvQBZOXHB+IaThekuZr1ieo7gpabRm+Am0AepkePZpw8IB
1aiSZaedMRHUbhX4pNDvc+cu465tLeyCrecs7OU3pX9guw2+n8oPCPJoX/Uf5lpx
f7uZmI1Qv+To9c8wapJGbiJpx8a1gFry5k8lbK5SpvsVbb7zUCdRl9NLrSK6szsW
us4fdLok0j0GarsJeC3Na5kKdvGHI4IFM+EK8eVhhKtLQluQOObZlkuluVo6ZrUO
T+/zucWpDo/xxrR6JIgXNRggJXvD+Y3/5G7tQ8LbHwTJmliL5/00TxshWqUuLRPK
gC9LsATjpZRwfH3msRHlFAN1MhGV7lplIv4DOirYB7XPdjjWRvNkbNgdHptIdLoL
Qcbj7xNR338q/wD1Zc8vwRKLloQRp3t5OR4sDUwfqRYDpRGSRMSsIg4TMcC1kI12
aFDapndf00FlxZTyT+3a/mrh2qv4u0uqeVAxdGUcqX35SJNqkKy4oN6WhpvmsP5f
+M+QWS+pC37M6xx6+0J1gmOMfovBeThtZBhO5e7tDPTkpuorb8NgXOQn1rRE3qkm
wfHWXxbP4t1H/o8Hy3SRGHb2sDfk2mVFl56VFFWK1sNtoOO81rAyGlS7fHGnlIU9
8EYGgCe7Qc/4718zKcLLrZ6eio4f+k1yZ41Qm/pA1rikIqL032dKvQhM9NoteObM
HQZbY5VABccfnzjxUeywsvLYHKnIMzBQMsSiuTtcpBbNpk2aYz40OMjA6NRy9Xk9
eV1RszX8DwgtVDIFfAMMkSEzZSCWTONGQ19GTkOHaOBDq/f7ToN6KvHoSZgpSpJq
58N1Waktct/DYXbZC6fZTWp79LrPTRBjaP6epFrF6N1RPngUC0XBP0yatYtQZSBP
rEgqN7Iaa3BiHIc2QX8f+yQUhE/WX/+yIS08TZDAV6NmyG8FhoK2KZUTzadCsd6X
iICyxO2WcVNiCCIEhFwUoHTPYQgQagk+XW/sRNEwuU+jcUvesg2LG7sCjEvZwzfX
SXduDP1oosa6Sn+2NLEZNwTjAqtnWG/kw/0/2aP4HS/aLeFmVPYMsNTXCmA0Zs60
F7mVV+9+cL08QSaZ31hXUMHdC13FjMyXa6hzD1GmOJpeBDJjTnqDcwD/eceWmJiP
YcAb0tULDPZ1IFkXgYosBcYP7sSlvER3V5ZGRDe+g/4oIDUpZIX3o4X1VJqY9hTP
JFSCPYiZ0H8v6JYeGcrFdrLdsUhsY57xJ7FxlycWUJysiO9HH0RRm46qoqdlJYsD
4yjIsHds95ssLAGm82tLE5RtZtUY4Tveim7lxhtSehoQv+8IP1QbDwNl6gngV6PT
0/i7tjz9JsBToH9GABc7E8A1SnPWVnXLyNrVXaX6eQnDkjDqVm/4nVxQ44mW91Uw
BlLyWXdNrvLwaXTz3z4hotmucVM/GERN/TNVDH2L7WR3OThblii53pafiVN2AvGE
m1mUdBY3mnZreLiIVO3d/DZCha/dJ8SW7z14/XK26/oBCIA1za+Iwg75zdRMvwIc
ecwBSUPXdA847PXzL8AMpKeI3YLoFbX6vdDk8o7gknN4Yt9hyNbj8lDAVpQKomFU
p8ejGFvfHGtZtPyHnSnIj7qdKze5kFh8OBxkIF0FHTYkHf7XIJhZNVMZheNm7sT9
TT+hAWk+uaYrk985XxVvreGyErQ5fcZVDsRMEcuznRXBH7Gr34JGAFFqvXTVrmGH
Xh2gO6poqwPk1aHPGWEAf1ZLCF6HqQXRXMOFMmKPLKPfvWZst370oXTEHfbxNson
b+WwhVEetIcz0z0PEvpoSuc0feYXBMYwD46vb4x+RgxHgifioexcNi83YYlvQ21L
D4Xb1xcRwuL9+jIILYuazB4YaQXheLzGu2nkKQukuHYxW9Csr9oBRbSqY7ovSyAv
j9PQD5kGOXBkERHk8iGJlSNaOVs2oEd7IOgrkvByuQZmY5pT8ANEY/Ghcror8VkX
g/nC8xUn3z94Oe8glWPjvGV85E1tU0bwqt6Ve18iv3dTfo34RQcszz3yvSR+YmM8
JiPriV2qU0TWTKemxp/x4ykeSqlBsAlzvw/ek0bciGLNjt8nSkYui3PuSAIQNZf7
Y3h9ZJCv+aYG9mKRw4LzKAfTriaioVQ8S3i/wYl/80s11Iyn/+KPALwwa3t8RgH4
1/GH2biCyARb1F2pGXHFdOhailmcaVqUFBK5N8KYmwWn2+QhwS1DHdSQp/NPcD2U
EQDDLUGVeXul89LhMM3+peyn+vy02nF34e4WBTtaqLkbUtu/r6AcxTBR+HW6M8SZ
AUYjj58wNYV50UeBYiJ6hEK0Ex3gjkp38SRAZQVgwzUgLOHsbz3lxWUb7e4rEvUg
qzBoFLfxbXPVXA0eY5+6VazD/a5HGjD0fSVFl5dYjs2o5eh6+oyxAwt7TfvbvTWb
VO3eNyUgooJAzsCI2Alu6em9tIIHS+uPmA4BJGyAQBGAmVVhUfIxhaAaRM7404BK
mbGWEGyP43nARBrnwGVLZ1egdGMosjxqBy/9Ab5TNHlWhsRRtJERZJQSHN+qd0dR
RGkjGcKXtn2KXUJ0Z5ysYSspE4K+WSNXHWgVAE5DC3CEzRI9qNp3pYbGHa06aUP1
HOWRf5KcUWQRoJZFzmRMvhySQch/xhsoEdCllHM044FTKvS12tfyZGuhLWTxzcHL
P6mSpL6dlslfUnNUv91A72++4Nksxi45rMJGtHBJdLUoOcckof9dkRVrzKReweYi
M5fUKLndCvRt9bYyuy7VREk1u50PlWPznupu2Xd+Y70eWUIHTXfdqtYaHXiogrkM
hi2GiyxXthOq71wT+2gS7eWzgk4KmkSna0Df+LfApMTWGPylVaIllV9WdmVKDtLD
pmRE+5w2g1+FDPvYWhsRVzKrq26+sS/vfotAMTF9i+JsVvDVepeOMrU2tGnEGfdG
J2EzbBOaOXzADctG3U15GBu9xV5aKWYRbbvTHc9zhI6X+K9cRpp7Jji/Z+U4Nc4Y
V5xo5NsMOsRSO7HGnbZ8ISg4OETkjwZSxb+gWWsM0vzWIDMxmUS1pNdyAKyFwgHJ
HrZOQQnx1hJDAmHiS5unlQS7fq9DhVeIsXo+mys3svlIuQs0zE65rn0vlMtoM6vj
x5BpFWr1+AngQwXcc9J+hJKrn24RJvUTLg3kU9fIwi9fqXVBr7CNd/QqjDenIeLz
MAZHwgj7Ggd7JS6DSiXYDyxcRZk2f14zBQT66AmqWtSJx+qcJziyi+wdKxv9Fvyk
21DuCOedkS3ecbuB8v9u3qEfcqfarLN4Cpr6ML1/FOrQsD0RUL0/xjKOAMP9FGyc
NX/eYnJafD7nnnTnOLlVKsh/ECNNemSRQULCAfq3t/RTAHKic19azkS+f8u+HuA8
0PBApHvN7A+O6rjTnIikFhAjlQ0RFgX/Frl1DCT1Vocqp/Z6vhUJKHnxhuSpkBs9
tEvIqZB3soLNkCLFjlos+n9FfAiSu87CqW6D4LRfSAHSPvkIbVsRdHAVKxjRxFkX
zngB2J4SwW0aySzPYcZ/xDcAhLJcjltzOk9M5pp3KkGIELaph1DssUGLBpWrego7
HMS8J2veZnoE/kAQc97TIPVQyT0v4LnbJsFs3dIg8/Fgv2x1c4xQywKUv8nYrHXQ
vsXFdSd4MuJlkiFR1+8IchHERTJIIuy6QwXhez3XZYuCpY/6Vju3LhRw6Fd5Fl6h
oLz3YYny0x9FwXfaIQxzNSDfoy7tz6OjMIjhWmYJLMY7wuSmXMHEHc5Ib08Y1JUz
p4Tn2srCB6tOykMznmksf8Qt2hueCvE73Mdvf+boyvBKSi469Lb5k1RtOsdmJoOO
eAuBqKYdmRpgnD/sQzqjxkfjsmABRgSav1NxUkHTrv06XNoPLHQJ4UGWyRZ3ReoB
d0jskWCZOpfoWXUbQx4txh8vwoV++s/um2k8AZEG8FiMQEsjI6iZK7/KiU1KHCpH
xpYkTtSGj2jXX5ChwDjLohjMKMlHgS4p00LfcBsOQU7fiVHF0yNd2V2NvKPyOKfD
lq6d/yuCxA0HClgMa+TfJDmD0Xf54TbQi3xGDEh/NaxhVMZMCwA4/bidKgw2r6x7
8BONnXmvR1q3ye04w2zXUmoOVVn5KOuLJVINvtiTrAQg65oK32m6lLyKqIUAA3XR
l8vFHwnLXI9fd42tUkt3mwBjrXK/ucVcLhR/UUmotJGf2lIsb+2jJl3ohRN0cquk
El96xipGcj6hMr3puzhAYdrhYyi6aenxJyf4SGGSx2a7w5QxnHgezSWP2Nyiyhol
l6LIH/nyX8oiDLLQ0B5xIAIAfmiv7xQZ1fZoG92KWQydRHo82znawIg78wkMt4le
MODvb6w+XtynRq/KQuE6XrS+nvRifZ0rRKt67z42KOT+CigMK0+janNZMrGnpdsr
VQvNeLbynagx2xO3rbsZjKoxQBuYYxU7Ij+FPVSD8oVJ/WLY8phdn9yDQpgfHYUP
nZUv2jtkudgXJpJibe33tBfQm3T0KUwu4reoVpNO8bBIOPKveJTcj1LE8A0yG64H
/PzBuohb+ooxFUHAKUezcoHwY8yIwc4GGfNjmrz+JjbynrDj2Lw/PKPoc1P8hR2O
tM5XMfixCYHeAX3eYCJwFI/lYtEeviAsNZxT9EjZuWv4Aep6Rk0Sf8mRvenma6d4
2tixjgBd/++qTMmiCfoN9T8+m3jX0EM7jQm5e5rezkwTWdti+jwhWURHYJyM2fGn
CGW4NPKzcQYXCYwM2F7qaOc5R6jKfpUFmQF8/VXWjnrZxs3Ma4VWx6kMyVTBd3aZ
fTufmBOm3f74L9qqfgH13bHVORLFeQZVY6x6/zISl2mHt8t+CSx6wyaLkMRepPok
1wQBZbiWE/2Z5KzzQIfIfZfRsLmhmNPa0kv7cFYRrDCJmM9gr8sN2gaDIFYpSAY8
H52uw/979hsCAYwd2HaFIps9ZiSltdREqUTn1jStyVD8TsRWRjDpecQe0phwaOPQ
c3nv1hLmaMSqEHrBsmis7ZAOW2iMZS0TpdhWGlT00fcrdBvuMOm9QsLKz+NXK08D
y9UOLeNTNIzYaR2i2OOkKw6KMJo5fCho4S8xiKLfamhNiImdWumlYymoyDaJTzr/
vOpXtmn6GNu01E9jNsW/dIhzmwerpv0Nsc4MsqhxkTwAub8duiT7ATEGt9v5BXZo
plFpRG3MRe4z9kZdKey8zgmcxDRXJeyecqnurUUyxAdz5X8UinulzxcZLIDQKybU
IFv0vS3JD/2iMrdAbMAEifre2Z0rqSZHtQIgX3BPzzOGgi1wOenrdef0CMVUjZdq
rHCyY71YTOOdC4qjJyUtnPlfWUJuu7IiynYJKNNloUe2mp5gnyQSiX2JvvtJu3MF
Oihxv0KwM/NGxHGIecGzQCMb/KBuvwZYbJYVATHkflb2Xmv5yI2rZyEoP2x7k8t5
zkIfLtoQVHvokK3BPbVv36wC2Xc1Qq8G67hl65bI3mXJ/4R0so7jjocSBrPQPFDQ
rE8PugSjBRF9qORH+x2CejC3pNZw51WFK/ZltpRCJfJM8w5ZVnDzJu+pesgKMecg
BPPeW6ZKzwafkPIeRba5aeQMEL/JqZ/rntio2jOFXXW9HQeekciUXgJzyFuyGIgv
tCm9fZib4mC6wJAIrLUCMDEpUG24cFvh3Axh/2ByIVoU9jfOcXChD0h6JGutaJPa
1GQc+YNJQo2GwuXTdP7kkm5EeMB/5bWyuX1rBnrb0L2PCifESc+Od4OoSO7kJp41
oQAUPZ+Mri6Otjx08mTK5aWcZoovHrSwzLUNV6bzxahlhvxhmPGfBbIKhiJl1d0p
5Df2yXDOvp+UW60JXq2oSqz/iKabLkUNM6l5Ot/lB7JTA3ubW9O5ObmlJX7Tme1J
utauLjLyxN6kX2hI1eWajZog8jFymSVI8/Bu1z8OPeQkiZIDRY/x5LAzdZQzJIyo
iAfsiSvhv41zLHxJZ1rUEjK33/dje1iIgvIkqtEuhgZskmIfMVJy1mL4i2moYhTy
m7WbNoj20rHXwynTRRhF7mh9/DlBXpFiCCfgdNolgMjYVTypD9Gr1zE4bzY7wi1b
lCoQ6vfyOXso4k+NMYcQgw26qF9z/NmOb9So3cMaOYeK4zQSroZlJ0QrJbRzGMcG
IjouxWMRXrM99CclQtGL+/VjzT6+MjpBMJL/3Q1f0K+YcNUT6lmhgIHVA+M5nGWT
YvL04co3dGaMsZWCPb6sCozdzIAZnrE+tfQI8pdOm81T1Nh7BnjIvRgL8T9HmuWR
gDSeWCo2DzZzLeCqK6LDsR9btmvi72IyCmWlWChvnyTXRSEQ4FY9ysiWWj9xwb8B
0DdyXANDThoPzWArkCcYAQcdKIeMvb/CZuVFxYwW8NV7wCVNFV54NkFKfak++hp/
rHbLN8iY/XWATouGYDMpeVOkDqz3qyGrUeEuPhNZwfJwTinjXEe2D4f7r1o5r8es
lWIWkEwFHbeStPvK+dNBg0iyeBz830Qm9AGMj1lgKmXZmt6fgBCyfYF6qlSg9nfX
tH/HL5rjLE+ZnVu2vhAZZBwNHphbR6L/gKU7OIleZZe7rwm7CEXOIXSWf/Q9+UgZ
tC+FwbNXH498x7DeQnNUEGDhVYtC9vtDyqZk9k8TUdZCJIz2wx15EjYOHqPb8mNG
vQ9rlNo44Z9x9k8NHnRNSpI6uMEh2B+nk1HZ26+v1ItqMKgXH0RRG10pwogoqQeK
fumVFMfuSw/xymdx0+VzCuVzDXMcXj4M5/IyOytXf1qAdToeB1OR+6AEec9Lb9de
keIamPjaPODMKTvLSuIzfzat2b97oSv8/HiZFDNwvRCE0PllgUXO9IBZc5YN6Z2h
y/oMObymLdVcSuGdWjMTYriMaC6rPBWy9zmkEAG34cevGaOrM5tKS4eUt35tArSn
SowtTpS7MkGi0ELmTHypc+xUy3Qi3KOHdwH+XhN4lpmW79BJ7odqEv+d7MKgwDGd
GUatVYif/h6X4+2rExyJl6mZ1HLAgJtw9bKYES7py6yx88tnpaSoStSyRqH0Jt7u
/fyR38h+do4X7wuNSGdrHr18WYVwsCmAJD59KOpsxdd4eGViTiV6FVibypTxiFEA
eSEG5o0QAXXUTd4cSFkugTYwE9yM43w/i9v9pEubok8Fdd5DAPfjF4gY3oJWk4Zw
KHB7WAWjYyqsKNWATUmPhscGzNUmutSg7Zz5QUnHI95/Z4TmHe7eS5LinnLZIFS0
FhxlhKaSgm4zasrCwZsCPNBJDJIOA3afpeCTmUfWpwCsqwFev45J3GWKe9nyU1fK
RM87McWiPKek6OBZAbDMO1yZPLJm+BkBjxMtyeNLQVFkG7r67r9yPwvaWWL+1TCj
u/2dRbO2HpoSkpx5r6Sc9Juvw/3MRGipFTpOizugEhEFh9ywBbNY1bmOd3/t9I3Q
9yT3NTeVcOug4Hnmicpdo/uV9ukvKANGucm3TCt/GDV20q3xi45vYVeSBzSDTRXC
fAR9b862RUIXh89W0kqMtn2LF66GsqZ1gPcM09uTdLE32igNjzS5lU5180fMykhH
nRCCqDw8+UDB9nFiZSAyiRTRLII7N//PeGt7GvxAN0A2fFJotteHx51gL94F51kU
Fur0SF6lVQdBerMzXoQBtogFeIv9lqGAyLb2ZLeRqjTXX0Qc5+lHT4vbLwcSg3LS
EfKGI68EWabNuaB1NXe6OVR64yb1bXALnQir5R8GFoH1Fpm98TqWGsSa46Gf6aZW
QsedbNXhXQ/H7tTek+gLs13s+pUroYk5+w3LRXQna4WuWNBw6UcyPeCDrEZ6j0Bh
E/oYUzWo9+a1vU+ACkSekCHIzHqc6N5Bta2tDQTMTsd204fnUjIftNCG53Kv4SnS
dgQo4dkSfkIkyuwXvQ/5kXQZjCjPA21/kzX0gx9bbX86apVM/v5Wufs4uMXm/83C
uhvtQwsEZB2jMoEwzkB/32iW4sf3TpwaGBqyVOIVeUSZvxHVYwo/iwZ/XUyi+lB1
iL/w+e5ej8wqodo9S1003GaDLBMWXRpap7j5AYwL8GZx2K7RwjJoT1IL8eGC6r2K
LbB8soLFsWIsHrT3fPgUhphSNuRBM3bS5s1S50EsZIw/jNAR0l3XMqb5ddWC2uJy
KpiSOU2v/ZYKd+tViMh1shfXfgZuINhHZ2Blst5JNwakMVkl2VvZoznxTHR+ZglE
CSDPA7Hssc15HzFUFtMh2eSQDcLARsPPALMO2uw2qLPWq7ZPHjsP7DGraJzB1CSr
THqFCvNzJt43/IzpHWGFkYxQTIvHO8i2hAAet4ruNbeN7bGkaQ8AQWBmNOS98Rw/
TILT2xWvuMhbMVzwXbqVVjviR14few+Y8zffZPc58LXZFhDSbliqzOZMboTRcOfU
YuXkSGaaVtW2VIaElbGbrOl2Vm5dxE5zA5URoN71I7uGa5EEDaX3ef0YVziIZDdL
S5dabks6HeZgqGaEiB0nVJQjqK6Y+dfKQO3R85tTYtzEL3KFmf388Ecm5ijXr4wO
nSU/hYokYA3j7r2um9hxjxPIpLA0B5uqTmVNnzdrNNWHKAMt7T4X1mSGXZlw7Mbs
aP+h/5XPSeo247SfJ2zhWowC1gTxgKQYLbu2xcMxwZsxs2q121yjoxgiaPxRLOcA
sSbv35gP/8fGiabPWX3qYLMerPeBvclEcRue6W7f6o9MGX1Dl3i9AudBNnKC8n7m
JWQpQxUjMZeWySi5mEf41XEzYTgNAqCH8dGU8eSmJ/Fm30NWEgo/iY3ojmo1OGRJ
mRx54UiA07nTgIXB3LYn4soZwN6noOeJQzc8PH4Z27jn963+gaL04U70ULguaI3o
TdKOwqvtMpmy9Fl92jP2ap3FQXbmVqse/drchLgVrHZaTfXCZFLwUG63L6eXEV37
tuT7e0xnfLvxg2SKDIcBX3cIzUqnFe/umlYFWDgie7DERY0k9ROnZzt+0rHqjuEr
dTnL0dbo1yvvR7Bg4Ba02ZlYD566pKztqot8KjRvueNHq7SJYiCYMeX66T7Xl6Eg
evfkUDMYl5dhlHjLy+BTSu0fSoB4BdkC1agKrwv9OzJAJAw3wIRmqhS7ZQ9k/xMX
HYVToKLIB0/EO1JSeHGoWODpQZodZTfBJXcBCfu6WUzexE7iy0Bx/tAus+wSUiVw
CcrY933Pl7+Ywdk9yNGbk/5xH9dDFFO6Rn8GtTVr0LCarobnDcX9UcRVAHft/d7P
JUCjB4mZOaUY65AEjHsRqm0N+UCc2JHCXBsOAz1vSNW/ype+9Cab8XYH/6tio6v+
1i7Fzl7D4PnR3qdJYYNgKNBvn7UCd5UgTHS2tNKc15g21S9/crk3xgnqwLqFdNo6
bmQxyEx359tB11uMXEZYymMTxzmHu7unf4qvYx1Z7yW6aHZYlU9UxAn/OMmcQsrY
h1+mOe4Vt3JDmqBOK+2TZFyK/tToTHs/NdoWbpQH/ll375eL7WV4yH9zRHiMd4QG
nRAMpLJN5cHXcVfSvr1sthz9vAwBTbD0X2bv6xyjDF3pWDvicd3WOsyuV0h/v+7v
ePnTpzQkvW6kZ9ko2GeoY1+DsO2eIn4gtaheIhB64AcB9G8/mH5yCwMzzf6JYYjd
OYcJ9B7ttK4olHEZ3BCLkhQS6MtX9PPEeP22Dev/jFnMNmEl/658YnZGJzyLuYvI
xdhI53axKcDeINBTQrK19UZ+O5JGww8R/4eywMNX0TCqwVm7O0C9ZTnl1HAb4QWW
xSS5vY8r44TZfDmCg8kHXPS5U7zMuKNcu6Z6r+S0NyXfAz6IIx0wnx2+Rvwh27z3
tKB0bUMp3o8s4wVu/ygjB6Z0nH02qu+En8S17pjbTKyHvUzFuND86t8AeI7bOvk3
1/3IJ9Vf0ojbmgF/fOochBHS7CY5Eokx4EcLych8MWwGz7nmPEyZ2TOK1Z0YP3vz
va9GRKyiClBvG4mzH4TK7WDKc8/l81Vefowxa/j4o0arlU/bPXGGaqFlw+jnsJgP
8bsh8Vrkoay/bNhbjmhCSgQJ2VTzBfT0KUKe+9/YPVrAySu2QmVCmPyFVm1/ka3G
ohLsw1U7K+msYg5PJNZ8eZpoqJ2IPYtNCa44EdDXwiZnGNLPxAk0ZOWaeR37sFjJ
g1iio5FMxhJK247MFdALlhfUlCm+PO8i0ntWP5dMyDQd9Mnzx4o+MUfscXCCBll4
RreKLe1nOWoK2O5/s+f/yttWASCL63ZxvPc7zGWK1jhBUmSOCJv0YtK3N7yLkbIC
4TJ7iFskXVBrFCzyNhuC3Jp7YGEW8ryelUnNUbpVICb6xktVqax8ebOa+WXVFGOL
ctomycUC8/8tG7bxWyWZY2+LDpSK0Y07ztgZ+0NDgRvPZtiPGBR/TxZG9pBPS2xJ
1YvA2nnpEqyPLfXKsdMtBLtKeQ+Q/wts96uMMiDcss5WKW4+A4vpO+aqVvvYViNG
4lWdoqL4F/Xg3Emlc5Ee2u1I2DjGTxurkGt+uQ/NjfsB1klX61x4s1nR2rgSt4V7
C8loHwj4ZsS3USKGAdzsM5c14cnHmrvf3EezreWPvhn45qqrHNes0X26wo/T6vVN
tWkoBU+tcLmyoqgve3GcvMxhzJaADeImRe8LOCzSGxIEPcWhyD+EZdsjuav5doul
H4s3tPm6lGCD0INDAIGHyZtFpkQDdTiK34rKtJfsbxHza9za7kOugtS0yN1Hx7k7
oTJf7v2y+j5/N4DcJ7xrkrYPPLJ7yD7xWvi5uDQuw1C5TWkl5vgbdogUZki0IONU
xN+RGMiJ7a71oHxXQOY7CJqa2Nfte7GqkUovjnCwjARm2RAGTNFrL2m6HgprVIr6
7ejnhpNyEEv/OTnox4vAGPpBk+SiFE5qoiD2pfg/E75AdimisS4hDtfdNltZ/ptZ
qZBtLd2itLiCDRUTRz0aZ8T0dNU1SqvIgjBInMeJ0mPgY/danLucSX8tugZSIskL
I1o0zhVfrF8gSMmHqLstoRVbXRyRwMyAIESZGPbZDg8iXKtiLeXGFf5noiXxNZtF
zxm3q4ZVh66ag22xpOY8cXpStwOIjPSOoBy/z9ERofXixD/BJjVUwueVohkKOtC7
WOHm96kDdM10YjgFq8HrZ062QayM2aULlxBlSt//9Ra63QqIijgwJ0HpkWGviXfX
LN0ozIfGDXK8CfbYwCky3gvuxyadWLeDo6pCaZ4ljpQOAmd9zsmQupjmQa3QjMkJ
VW1gE3avkLZnD/J5IsK499b5cQCdouujZVE2O5vXkxu1Wno3GdNOQmILnX/iX90v
U5saWUXGlDPQz4vfTOfqyn6R0TOXOfci2KwjE3aMONo4zH+A4/Lrog0KF1zE6TvQ
uPMUjN/RKaBETv0uM7wEWJTug8ACq0Fq1YRWJ09MY0Xgw12aIsBBmZJB4/UF2ldE
mbscJYA/58tIkOWoKadxtn5NLL08lMDKUIR9u2D6x0MS7OsPwliGPz2uW0zGCesO
Pw13pgug8xW+R9En0Z8Egal63iWVFsTAUFTyjHMO9+OalzMSNQWMqDXe/ek/b7sV
0dPmTx6OX/1+1S4zyOQT26mcnCgGhJWsXseXmGWBTzy/EdweJzAao7s2XoQxxua1
jvKDqCXZa8tJ4ILaYhHISiXjNCQWhVvhh0k5qtMjc7SVNKOhYbNjDQwgmV3s73V2
SuPd7fVMV6uy62npbeiTfxpXE3Nv+JF46dxyTRtnjjk/sUuBrxItlDRcKGt2fo9h
af0GDxhMjnbzS8Be51xumDmwL4D2uHreR32WSeYcVjB7fUcH00jhi4QlSA2X0efJ
pZWauGiV9UFVBcjDU+RCvEKm00bx4Wl7hssDhgP7Az2vAw3RzyBldxg5nJ2Hkevr
VFXZx/zRhnAGRQmOHCvDJPa8HagKlzBCVqgWEhBsgJb6jDH2LNveOKllrqxouGrI
YNumJgCoF6y3ihrnKMsN4hwZM1cq5BaEjDh7jW4bPszvlvGn2mnA1gzKQkBuiSP8
KnvY2+KOAyphigLa26FMDXvFJ8INcL1JK9p+D8xrWhxLz/uIOvGaVgs0IWYhSLG8
8O/Q7bVhkPsux7dlj/ZyCLEEk2M8lbdoOJgyOTJkUpX1L/Vou16834YjMawivKox
vAU8eK7I22ALaxBTbAkl5u/4nJN6Az67I4m8o92ig5+CwRF7nAqFVdBTTTH7P49G
b79Kp9PQRt0xdazQpOzwjyQ1iBmrOAVkExWlp72GABM1uIeRGyDygEubKKXToSL2
dUEVsCE3WcLUswGOd6v1zPVwkhuZtuS7wTLF9/t5B5ybkER0dkEDllBw78ijFmXJ
UB4PTasONescb2E+oCSoaV3MCGseQM0mA4IZLGZ+t8u2JacKvxB5vTIVi9/tVHTU
2qzj56bIAjUsxdIDeuh0uF5QwMH5u2Pqjl+JVlJqsZnJX01VUKngE5SoI/O0hV/0
+kGYcnigyygZtOgpPd8fwzKjg+tlB5uheuMsslYccWhqhcmqKCUfL79BJpfz4m7D
Mr8zHQg0ZAk7fAmJi2AGsOHQbgUgZ+lrq3LOsmTRGPT5IsjV9JmvIZ7l9Adhykdo
KCRofcHoWX2rl8Fsqw8LomxYB6MkLMOj54kPkJbYQAm1dJ5dIt3S6esnTpYy+CfI
ET3qIKbPXaCAF/RDsWgjnhYQpHf8e7hM62Ckbb/wtFUkOaOuOOnbelph+hPbD7Ox
wOs0VVYr1lt+ylWIXis7RCl350DiGX31mMWslUyxEZ1AxYdTC1+jAz79JiFMykEu
iUNEBRji/a0scjXRzuvNUHWABS+9jbBmZQFMuhQyCvN36M8zjXno9+K+HCwVNyzr
3YLyG4gUibXT77nkLNjCXcpTJoEERRiC9J941Xz+ndcAUFeI/V61/K2FEK3VbiYL
TZug4kfZA0XWMFJo2015uzyrJVjEVxItDQwwNJefHxwUqCnzTeSu2/rMnyQ3iziW
GfFUmZSudrFXGBvt8855INHOGPwstm1vLenFj/vn0rMq4+fGObGIGE8D8x0pzoqH
wDcWOJpHIZ5SmwkoOipDaPPujuELGTnX569OlyNTdXY7biBlDQRw5E0ondytN/Hg
m/4wycbvIX4DkZQgaYpoL38RCYgh0TIwitlTerVYys3Y6dqbi03hMxcIG6OLeSdC
E5yl2NkMtYbkzAjBJZsS04Q8yXrzRSiuZuEYLS9PrzgRH9dqr2yZNWe38Al75DZZ
EMG5QogKq6vI4y+MMoiLDeUgnL9VzxxD2xDgthV3sjJeJXGRnqqxOJisFwiUaKdz
Vxyb/se/zD6UG4LgWSo6MGqU+c+DhRKi8fRc+fKYY3lx4DDQa16duxNuI+C1l1Rm
uXg05VbepwmKvx5k8pFxMTzBo04Rish09ztvIwxYHpfZxCvTFbY4VOzamg4Dx8dm
FPAZCHdFanD+tVPpeL4ax4aqsELWGOz6bRbWRAxcva7WelYekURod/NCkmt8dH1V
q7ES85SCAJZNVktVe2kHXN6UTd2dg5ljMr8NuTUqZ+1L2byJUpH7YZPJanpBIHAj
dmj2xce2+B4DuejzkN5qB9/Nx8viIOYTJ+E7GdXm0+VjUT0Pl5v+nKNxzJHSPvf9
QfgCgL0DKUU58OnfAOCY/EdDgg4rweOQICfKGry0MfW9PR2eLBxDCnyq6ITp1vui
hY7ppvW3MySLwFkaP5BrZjIoym9YNkuQnG2ir0TPT/88rPuQRKaOvUAUx4CsQGFo
ZQubFNblq94utfHhXfj/7sz09HMNHlHj/RHMaai9sr7rlltfYhCjImZQi6CCJzDg
z57Km6HzI7pq3dL2xosz8sEhcVU2f3I8GFAo5DMRyaTRaE83xFqnvSw6BKAgXF7L
5NPlj8wdN9TkCGssj8QwB5SlNjFN358S2QBSHiGeCEmZhd23np70nMjQp8biQ8jr
a/HrjvSdkT2Kx/IE6soIyE9/RmR0ay8i+FUZqUNaYIIIcmEDExNGmj1fNeiI8lQO
v5j8jLNt+qQ2qeYjt66aoDsSuD2/5q+CoyugswaTatbr9VrsjTSVHVuFgN5HstI7
gOEm/UA2/MtSR6uyK9SpZa6Ko9PaoI/6RWBQHARi4ijKYUxieGZCExCG+E0e9OBm
92ZqwFiNPvagMXKN1tk7BRaE98xiZuyEHB9dHiSpOjdSsrHkItw5LgWL9ZKWtV3Y
u6g/twwe8DAOFJKPps87+9PBT6L3sW2bdxPYaAl0nJJby5f+Jgz7dLx2Huz/CL1m
bvfOBmveQ1/LVVgxMddWmSz9h45R7Hc1DxZilRW0T6GgQX+2ocI2YfFUkt7GtZTn
LtLIkMOevxG4voipPjTMFqjBE3cwrSXzhyhCfrjDvAz+/EaHwx0t4jHfZICixpy7
KIHWdl08jwtFHQtZ9Kzd4ShVMGfTH+ikX3B1SioRrCbqxN0DJZR5CxJF68gAqCr4
qQkWbTpLCktCTaCXiG9ul7EO89gygwMvtpGucQFYCpL6c9yL130hAzn6N5nuT9jm
9GLhkoSL0Oq9Lm6VtEQ6JRBqjwMp0KFmwejohu63/iJ1Rp7glf+9b+LDd9QZuYFU
B257x+cxCPC1adY/6neXETcAPSxvnI7kt0iBCWcesGUuu53hmC9zP/ifO9LhnIbw
JXMHUP+p+aKy8fegAGzNiqRltI7N5BkR8EeoEZ5tpulU2sges/fr1q9B91d1zU2r
eNckIRWi6uANCIWdPXsoGsKe8yXly1SPvFyX0V9A0C6ZAUDv9bK/EjCFGszNLcZi
WgNQMTex9l39SmZmdkXx66bW6UhkajI55evGk+v2F+iZb8Rju4wRG2aVdI4U33Pi
/Muw6J5Fr2gAVNm8tBJiYx256BxitfLRfZbShCuN2ynY0vIk3v8PLdqgdthi9DE/
FeTSN5Y1zaLwfb/QaRQihURRk2vamkef0k8qU1U5wmpGTD8t1ErvstYXHEN296dV
zPkkEHzCZmSVuUAorI2wJQdqBN0k8Xdb/Vgh04aMoCP/+X7g5rKSP3lQl3u4vFgf
HpVlOAYHH2K17Q55N5jw7aC1Zz+b3ktO88Hz7uPVHHZWmY/hwpTju1UFpa6JEs+2
N9EfvHNJ2s1kd2CRRrpstDd/5PzL3DNCSw84AvGhbcObRZ2+5nooC2xPuAHDTTqV
Qjly4z/U5qziyyj/jQ+cUnLDxbbRh8npm3ceo0bw9USbKPBAmMrWXTAsoB1HGYtC
DJsTvBx86N1V5zFs6B7SZJJlSXqLEzBZgn7leR9PWM5JjE1/cB25ZtaoEmqJp/aN
r8LjMyyVokIQVywhdd4PC65mFGBc7pXiwWIY/8MfnG7PZ0NNMz3DRk7VXrJhsLkQ
2jvmMMYCiXe2qUGh20Pz3P6PRv0MXaLMEBm/mVAJtfx2ELhoqs18JYwP4ZEAXAnw
LYqmYGeU0Ye+MXW8zKD5MoVGPdVKNeV6RwoXgeORHOrQZJsgsSQdddf0qXi2YefN
KSI9IP0u/vIkH3CXpMsWAiMqKVSpTBqC4uyvfpB1itfndF6x1OePbfiOUEzaeCIV
igNPP+zYGAFMVdBLmjkfEH8SEqjaWS+RFI3ozn7t0kMM/1MA89juJc4wAzE6z5OC
JmY1+GnKgucayFFav7zFz3TR9TMGmd8uaXTa9ZO10lc151d1/iXPsCoYTv2JibCy
9vKj0DeHlujplhOdpg1+N++ALeD2/eMIQpYv0CW2zJRNWirtlDukkSyvHz3zPeKE
4vKSO9RArmFarCV+t00zcjx2DqygTmbCwlrzMMACptWLvnRe7EAT2tULtdUy1YDU
Ts+hAUb5PgD50p9oa9Eca2Myy5M8OTC7l7ZVU3MxmZeeMAQnTUH1BShboskRmvpU
5gjmFUZpDFrJobRJHn5R1SvQUSh9K8Y4GiylZm/GvXBbEL+OHVU+mqP+iBNnN8M/
N1D+DcSheP2TpYaNUnxXWrNaTJ2BLFrIX7BO395pAx9ncv40/c2rldDb091EC8A7
bnKzj3lGEOeDVTFwqf3pBkTerZZJv9EJjUiVPgIeJKL4SyebQPtjXjTzd1COfktV
h4FoEPwHfhuTDjGmf/OXXa4QFse7OCWKZpvk4y/GJGeqWi74g7QvDJ3/nAjQsxih
Z/+wFMQ1ihD9BO5caSdtybxc7nefkTSTP4ZNaMFgYTtD09IHwVUaTUmsDE4+N7a7
C08ghKnz3Xb/01mnNPiCh06NbijlUAMzIqkShH60yiegczmxNy218myj3KmXpb1w
8eJdmKsUJEuxscM1SdV0ePfq6oZEsQtvObmxjjN3FbkjH0lzWN2n2W392aPRFFhv
FJfKzwNBLIHCklh9G+cESQ4SdfUbwRidujPI+g7y2XZxffIUqlJq7UBLn5KE//Jo
S63uH+r5lMV+jvUFRIoPlX9q46/Oejh0/bEo6Hhrnj5jrkZL8SwphApPIOBg01ln
+PONOd3VEVQfhNJP8PbRaoYs70ia79Iyzzgfel3AY159JCeNT0mxl9we+SqlpeIY
iXkm5yDunIdQNiJaYfyovpQU4MT/AnnmmR2QCcaaJpnElD/GljWCTZvml9er7IxR
gvjQ3XB4ROTjxBwotR1O054zXfWf8LqVDks3v4ZA1B6IgVAevQUHtBF5aRKbn1Qx
agWHrVxBInQASFmkKAhsp9UmDoQdpRTsPHxalPu5TVMKyplyI99Vwjem1NDeh/WG
lmoT+WdM3tSMLPVDKzn0rY7Pc8IlmNZ0V7rH/GjQgRhKc92CJHxgVammIkNQl39s
IpV+lFoXnsVx0g0pODwlw15vWTmAmQkqV57YaQqLI/6JEcDHb7lwYUZSY1zwmXY+
NEVOxHGI5L8DHgrG5upflQGhxLCX8++8a43CgHyBOqiaoyUdV+VkriO4rMBU1QAs
XXls6aL8g36WzxtMSjPqFEcFrc8ppyPmMLj4apulT4wgdkRXBYp0aFiRlKSf343K
QYmZbzQYQxGZnk+G1yFfgkbzT2XiiEWq/g8hcMXqYMU2mb6QrZHVNYdscIFxInwF
mbthVJIHfNj1jZJhnJMSYHaxXg9FUsREkISb+JG9hrSxZkCB5TigiiRvybFQTQKx
a91+2eJgu038R4Dcr70trLf2RlDv0ZE09hd5MSrMxw3v4NJJQo32JXBcKjgIZhaD
CU0YLzazbW/Qytyv7+WXBnaanBWWQyNRsYDLwNhls9mAytQm2g3juj7grxoC5cQ9
+7eGmNyRTMBkLwdAzfGQgTocGVa9viwtEtk67AyvrmVjrqY3fkscG1RtWzDIvZJK
g/etmT1JHlqbb2Yz77MjFO9oIimlvQKYrcDgHBeuKV2ZTVu+5zG8SB1BnDj7Jeyo
OW6Ui34YK7db4/zV1oasoEk3wQtofoOeBMC3LFEi3HDw1g+/yhFdJn70rqw78MiF
B6MTtKlkZTx6qxfXJK6uorkfI1kUCxz8/hJQD/PpQXt+0Ya+aDcrGCaScSMNFNDb
YLI4Z6Eyyno4ah4rUB1S8+bRkAQ8b4l1TSUZKCrcVSEPZ5nyp0mSlAZ/UgigYJqu
9Al0eP71SRGI7OWTv8Knhg+aloWO1IEotVun0XE7ka9ifGy79O9oPTNxXBzXhslR
heh3GgSvVbtSYdLOG8m3slJu8AGuKDfSmkWlG+3Eyq/d1hUlcnRyH33e0vMi2LMn
Qh8VHAv+rYJR3VIfmAlfzBbyGq7hwn0h/tj5TWtLAgCg01rZc7AoueNYPGP6AanZ
E02KFFAVIa0cqeqk2h3hMOJzM7cqtTTP27W53sLExogAtALfO5XD6XuN90Vet0JE
SZA8evap8sVz3Z/foyclguDLxv7oixodTAYPFM5NKEtkxaGOq7/3hPV/Lc+xb2E6
A4kvRu4ynpGYVgfMF0LGs8c0HK0AXkjcyxf0eFJsDNgbCAkj49V9mAAtT7qd9+Is
fPrPBp2nq6KW5Nm8A4LBZySJQX06RGAMTmsPSDTjbGOONofDGcoUThk8nIrdIByj
Z1Z8zO2MFVVHWQtcwO5hdodzIhVd37445MhQ8e/w94wi6jr6ZaWU+wG7fPISyblw
3kGgdUsDI3Mg8eu7gHsNWoByCI6DyqCTsrWBFtYWqHt99q5kVUTRuy9wYF29zZHp
2VBD2uArjYl5aCy+ym5kcmUjy00LFgXfLX6nPGK3kTiexDOygne/r7Ah8fCdBKVg
r5sZC/cXJ6Hup8KiuPDRuPJwpxHTi5pys06uFcGosIwOvplIvKUiPQQPF2R9OKL4
ons+HQtYktDVH06Kk0JmW/Ewxr6FRQjH0OReKIbD/kHW1zn+TcToco4QNGaIsV/Z
DB3IN/eCwx8tgpz67YZn9JScPQ7cuDTjUv+Yw+fkG2LU8uGHNvzG31biI0CogPdS
VIoxKMd4y6WoXgL08I2DGU5sBhEZpdhfT3LMxclElaBhFxe92cLto1w/g4jqcRPZ
gtk4q7Wg1LAer1Jyx0ak5/sBNbV8tARSRw3H7CXT6cWLu6ITCKex7TxAc6mjyA2k
dTW2/1SXoB55WXS/kOkOphwUhms42P8hCXganqat94Dlqc4gOACY+MI3atTeVDmT
FZKRvQ4Yx0f8Gl204cB3ZP3FmKs2OYx+SEjmJQ3JJcp+ZcN/OYHovq/20nDwk4u1
akciewjyjBCPkLGbClFh0bpSJCeVIhs0NSrnYeqi0/gyCM3UHhmqpsXKXMa4u61t
c13cgL4rpwq7K/VRk8PcpzWVyslIbK73Hp+iaEve7TEJwJ7QiOltKu84/oOYQP2Z
ve7fXffL8g/Mw7Kq1CnMLLRhw8tJrmOwUSoZC2KX4lQrXKppzVYho/m3vZqalLd7
f4K/hV/2wqAGTVN6xTr5dewb6uyFzVlzli6wNthkguMvYH0lnWnNCyTL/ypIhWQ3
YLtXCd0coVj6MMOWaGWRB2YUo4/awSD6eSbi+Jp4PWqqtiNHRb6tDqLZxoQ9f3rX
7L5VBWkw2PdCylxfLgYLEkpqqCQ4ej6uz8VRtlVOhJJPDazewxZ8ys2K61KSUruc
nZZ5vF+BtWoahbZchdUBzrLLIY6nJociWlv7opbG5J4+PZSZLTh4kiE8Z8jkKzb9
dCXBti47WhE+iBr7P06dV+pTDlEP2vmcmAcEM37J764AITPtJq0HVyEj5bR9vjcu
ax7huRVy7JjI+0iIcgo/g97dbJhAWw9Yjmzii746LPfqZjmbWoEiik7MWB+4wgH3
lKPeYMd3OGTd3cpMRp7svBNafUNvnXlgBvHNWamsyan5lLJ0zFvmT1MYbm8w88zX
qQIhvgZf/4ah27CXVOdrdbeOiRyRVVKzARtqwq7kS2ZWJgH7W279mbK1P++xwgxQ
z3CQMufCiFcbos9FiOyeuSyQvZUHwLOOz6xi7tProIphCA/IF3U1BOx+rwHPh39E
CbVCPsy/Osw0tH1fStdYVDhGJ1Mm676voikVFEV7tb3CjFzMAR1rFZ3PheXJc5qU
wDcIuIHrKJAQyg3RMLjIa7WaY0bvVNupjGoM9IpxDLgesmTxGkHJ9K22ZgVVxVXz
oEu14SabTYjKjDMg73k5a8WrhRY8EFYAluD7Gj49NurrGkhj/wRYZG6Wo0L86BWA
draPi+2gJn5FPeZnU/+/P7SVSZKdFyP5yNGVuwyxXcGhsg/2SHyKHdMJr0rIiMdG
HpiSys2ewH3BxE6LclO5sxKj0C7L2st7tjk9QbKLa8sn71oADkjHybKcBm1EKuLT
Q4c5hcM5hf+Hn/tbHLjvZxU6Uh5pDnaWTii+OJVDLQBLCQ+5Q3dATOVMDDQ5cjid
jsfBlNichpVl+9JBENPLCblV0sQScHVXsLuWtgd2ev44mbrx4R/1tDi7n029YT3m
SmViT4bFJY1Y9vKTTxxuK/XM6mXy9EyfhQ3pusKs+lkKxbJ2yYec/NgU900RCrxk
K5J+nb2Aoby+x9BUrp8xroqz7MMZp+YbJMfjqIhL+ic08tP5HhJgxV1AMS2vw+Mm
n8xIRrY3dYNmDhAJ4MORJGZePDxuMCil7CVKhFtLvo28StqhS3oybaFnZ3P3WjJS
Zo2EaU3NrSFryi1BdcCZmQLz+xm4p9peUnO3VgSkoqCd3XlfCcWXEoWRbCuQO0Vi
hbhX9PXM1kV4oB2AELOpmlAhfOMMQJHvtk22SJom8P3KUUhJhJdvmjnazYeEsclk
Rq6IRa6noZVG1U7gwhMzCItOqF/5w3z8IHbQZwVG0LDvJCuTI4hwAB8gXV+WwTcD
6vATTcxkZBDvJs9bsQr1I7CXjjaiaR7hMvlomqLIEx9y+mj1JMoQTgon+Uul9ZYd
TSKsG1CmsTm5MZDOlnaR68fQrTcD6lHWVaQC04mRvBIh/e/Lxw2hZEZrxlNCXJIb
sV36ikMCixjiljwKqxP6WWFpLXKPJszS/ClT6hInqKSBmC0ieQweNSzoM2r3pAW8
x6j4u05jBm9pjA4qCvVoNneRh3dMGeupYCKm5sDjrA5RdtEzm8Z0TMiU8XahJAC2
tYm8Ts04HAPCRjSG9TJcjUzkWFNgH6Hk9mEyyO6vAh7vptORAtGzni7cgXPJo3fv
iWo+ZpBXlOzcjYDDbbCrwtMMk/vLXRHTsoSRboHmBQ8/BqIRMNxvDZ+qxjc6BkgD
p+CKetkuLCkHMwMlEyx4wjBFUzbZnzl0VXY2hcxz0fecJ7W1TNfwlKTaHhTkT3Tv
xUZSuvNgaWPMdXWTR/1fxErFwg2Kq0Vne1YogspEMgXOr8SyJ1wsXwttKm42BAii
Fr6yB1dvv3EZN9tzzuxAc17eaQq4oHAnSUziWcvaU/te1oBi2EbvI1qBL5kBv3e8
R1uXGIAM5ooASNc3HRkh/RzjoPkbe/LHBBJTKF9PJwFfPZHbT1alMzhfDF504kDW
zh4XEXqDWu9BrmpfAaIKChlmgfjdK+rEI7NMEUAzAN0IfWDvTamqQwp/R9CHjCqT
kjknTUGI8WdHIOQV/jKgEtmASxHlEU99FE1tgko39PIHVUB2Z+dUzgPn8eCB4Oak
w7fCuC6HpN7JC+UqxV2fS65Nz83RILXWkVKYnvH1wbFvVB8PaOI5SgW777SpGKGl
JFbaoF3vDNNdF3zAuiKFqlre29ltp6stof2vt/TEvMHha4HxYaRk0gAwNaYhSREQ
h4FAmnVkmTD0Q2ct+hHE/1FNsI1XQHfdOR7CR6Ll2Y/AgdSG6g4stuXFtqTRzSEK
Etltclhr1jSTaOtv5rrEy2fnqZA3fVrrMu2xZBIxY4pS1qk/9OmLMJhov6USBQz0
H6vUT2shAOCuOj5IBTy5/vyWMszcCoLrRXBaj/wQA5tScMU1TbzH3jwLKBTRXnWX
K+unrSQVz17btg3Gb9IZftVicCi39JaT4L13uiLc/2ThBOnMQaWUqSdLoXDi+y2H
ZnPFttC2HegtioqeTCVCxKHiPM4XtneKWQFk41QauoX9wPIyZJuehfwygfDQ8aSy
hgmf3AgGb4A7D08PGdN+3VCpAFEnksVKc7o1yz9MH4Vwm2U+1wh5OvG46kqTHb+1
iDeP+Sip8inLZyDyBnsWRMudvcUJQ9J5ezIdeTQ5Oqp8ZxsiX+tuWz8Kl0xCPY/C
FgrMmP6P+zFYbawoXetZ+SwYP98NVbrswNmJXvpJUD7V0yVU9ZmMUeejysJ2Myft
hBmUb4ematXp4GQULpgCRyq4/e/7YW8BP5ROldRhbkZyd4lgE3zVsWVEmBQS2wQr
PAucxEKb0nQnTIQLDp52+zz0fy9eRpwKj4y6kljQNwvUsMC9G6LPZo5qCXD92kj8
vcVFvu+Smr5x9bhazTeb/f8NE4WfMvKC/6ru3g5OPCUHuC7gAcoge/5UVKW+a1RP
ufXGMiwOoXBamjQl55dfx6CQWhCuoQpzPv1Srhvuv17qWhXEJdMzYEuNc+B6fFAu
9Snu6CF8XKXueTm38rYvdPeU3fi5lXgnE4nkaFXUXdHG5PQwpsdxWxyGQZvtRY16
4+HMU9ayLgMU44bqErzpxDzUSkrjmLwjCwpc6nP6lftGweKv/j5Ts2iA7hRdm9uD
g7dI0oK8Gd7DAGlT1Q+QeWEteNOtwOT5Z9D1E1MiUNyPXYZuNPK2HhDbTRbAi77Q
elZlWikV4us58ZzkI5yYc1V3+MriNqfH51KoNEMgklhzvX8/uxAYkkVPcKAv/dmE
wYeYwr+91eT9p7EWf1GEfBMvAPZezfUSo+rDyrgyy4kmiqkgmdrBm3ki0hnlbnX/
AGVgdScZ+ALX78NxEAuH7HJTlgICiMc17Dj5SY4kquCFYxbCYusHQOgHEq7y1mrQ
LtBm4H+eE4vgsDwa+nRFLOpiTv40QrjzpXPg722gmQdXSMx1N3brDHDA9AgXQJvg
Xyx+g20CpQGSO6Zl4zl19gXJlSEIf1888HbyDAPgDBtgOCzTfthKFWp+VhrMj6e8
HmB1//Lh91+tyWiz5/j0/2BCqnwTZZ7VkBQYW2LvcWNJvkuCsKgDjYtfEafQaxSx
TrVczCBn7sAEV6cA3gDlX7NxpzB9aaSOK1R9oX8huhHROXLXvYmbjGsWnVly1yhz
Njb5gu/k9ZqoOauGFpiETMakVfG4cynV8oI+bFoUugOGfeCcCJA+bzp/cyBF35pY
ujGozaBhGToOs5YuERWQoNxnLKfcRcaE8IcKDs07tyYDq6+G2DWLyGlLbs/ejhAS
M2vmCd+Yahk6TW39J/Jbocn25mDxw09GvClyoOG9fy6S9EXTpuDAPrFl9u3W2Mng
ecwvZw2eZjJ5uuapoLgHmx5Aap0qJsx3dJEbaExs4iZGZH0XO+Bw7jaXoZLw/E27
K8XP6nIjhWr99lHnVgW0NkNSe9GEc4LrSgT3woWvtd+7Hd2ykatEVqcagSxlM8bK
y/DdGuNR+BjlxPkcVxx7BOYnJUqbLfI6AmEaVrY0rrFKAhcDUE6VbZHoUjrv+Bpf
nhEicxdffpfFfUpRgcCwN28+RvcmonxpbcbDyGtEntBtNZf4Q7SlbtbWAzbeuMK0
tabzwT7nNmH+nq3Y1WcaHXfVaCNKVnIsF+TG2sj6TfpMj4JJtPUbe2borEmxtTp3
1HegOmSuzFz2aDzVRufT6lx1myj2jzAlFqE9JwXvbagpyazHoS0vXxd+1GkhFyPt
RENwbWwhHQk8x0ji626rk02itWC2A25VC+HzFbPznL7j1sxgCykK08rtg/+2NDjv
nx0LF0SdUBMFc3sg0JYS9PccV/zXpXk2HD1TrdQzyT644IrvQZropHQqOGYMAVzl
AjtYgHWL3SYTyepSVBir+cUuB68OLl3ZH6eCH57168s3kgYUYM+Bm8Gq483Uyoin
N3m30Wi20+ezNmiwvrPqCYIM5rjdWypYxy8+B12I7XbXXaVT4Wa7cSUfHeCuTJc1
IoCyKfiEyVhJIsleJHQC/81w2xWbhGRq7o97V6p3jnEAEE05JgeoWTKHn0TQhDBg
ulKU4R3AK2I6zRqkP7fmIYp6zAWP2f+gCBU2PdxN8AYCmZ5bL08tMGMD8nnK4YK4
RZKu/CvNe16HfCb1qhZaB6RQ8UbDxiHbwr200/YjsKnV1lFehKONC0LbrQY0o+Go
G5bScw/ZNN1RTfuPlPJdNXOvRm85r/n8cjHG+p2NeOUtS5vcle0yy0kp88tTP2DL
EJSHkK4zMd8eu7ghdZdJN6WD2imRV2XLMVA5RFK/6SuerAS7fReaT21cuTdaY9oi
uosbqFYVZXyYnQSpJhacHR1gKh7QG3LjG1WHnLq9pDWwnkoU64ij61xcaba5saBF
BtYY1OWIVSuuwnaMQ/iyGGATpXfndIWPQ56Cxm/oWBQV9zpB/YwNlCFFtdWW7Mnh
3Jp0SULmhcejaQOYbvPZpbNFLZOPVT4MQvjJWz+mEHxfNCH/eeYhXk/hj+5lMAc7
4SrrUykdUGNV2hX3Qq+5/9I0HrSoVXgQsD3PJeNQVN0BJWvJgXtaRa3+rQVUkYVg
TDUrGSweJAluis4J46Tlb4Zw2EmaQw7K5MRem1GsUN/50g8g0SVfJ/idz2n6OJJJ
ynJfMbBCqFjL3NK6lOPSvMC+AJSbpugaKhK9c1fgEyN1Pa2hCVUKmY/oSc97akCA
vj/At5lOL8bMabWxYqhwGZ5pmCe+ToHrkNBvfqeYqjrQkUToxkHttLYj27dHqVMu
d/AkouBk4rXZZ5a/kKx6Lx7MBD6r5djUWOSP0OO8sgrP9AkinRISXJVokF/LxGBB
t3nnO7vtA1KkFJOfpxfTUDa6TyXS+7xz/T03TEqQArRLEbMY0yYwDnJelIciBiqH
MYWj48UCYnwiqrcgYDhnuUeolzNHTzW50p96ulzUCj68pLr8emMSP10Gg0beCMfq
5eKPkC3R44mB4QS6NycTqBlUJ7F/VIBVXEliKtrHJ7O8AjBStAt8Xh3fiu3EnnGs
svVLZa/iIjWiaTqHXRixzpFjOZ86UHH5Pp8j2d41MpVNdzhsoaqr1Fq2OCr50Oy1
9LtCFHBHoNd4juf8/w78iMK/PYvqUKJQa2ryt9m6sy+SaXNDiIx/vWk3N+krxaaL
OVMkVXOYf6tLq/6sMP2I2nuMfVu6XoitLlWZpWrkYfwJUlXIc+e1PT9tqFdvB0S7
on6eAzw2AILzSmnIpB1AY9gDrhCpnMOFvkszk2gPwImQrnHXIdrzd9bW9+d5LkK2
OwgehXnbrcC5rT1guYEyhhBizyHATDkX7FqE8nyT77JtnpHfZOYiMerihD4pqzmb
PhQU9vcGuzV7ummGkoBMejQgJ73W4C21D7lG8s4Q9okjdfHeaJFtAvCV56EetTzS
4EukncskDR3uIgcM1u2JSpunIyZPWoTiVckJsbeRDvkvYKe1JYLToCFcU536W1U+
0sr3/JCg32OqGhqPC7rFLHSPXiZ6Q95M9+S946bAWVIPgJ9tLoEwaby7AnaPpSK8
05wwzOL517NL0/hN8vqZYXGUFsc3CgwdGpQs9wnDBdm/MsuwT4DRU7cJ30dmiLle
JVR6iLiNZyy+1UwtFTcRO3tcKzOJyBkuLTQ9bADGu4ZgrFbqtWcfNbkzxYX3BZbY
rThw/OPlH6TCBzARjP/uOOJHcAkw1nDiitMr4J4fnQGIUMH3rNIlYr4G7XWUE9gU
QOlzepHcjNyAaEvOUwzBOqeX7IZUkjWun2jj7xLMZrDqkPH/G4zdb/k54VHi/boh
656XjK6yUUYBcZp1qOxfsa2Pk5PbBle660nCswXsaZuf2mtu1r7oS9tFrPUBtcw3
obk/YbLculWVsfdZozucM1DPUsWZy2dxaZmyaNa6Pf4p76QhC/f/Xixy1MJWC22P
foZwUwV6APa7E3HrcSFhyTetw88t7m7Vbd6qs+P7YgWByZHHydM0zuKtoBuD7lQE
ssyVatqsbz8QMcV9ABwB7YdsXOSzNLZ0BTB42w3+CLGILLm0flUoTT8sUl15UM+i
tw2pF3LN5Rv8lGdqmnMNcEsCxrQubLSGN8ZhTQRcSQf5Mq81J3GSZRQ+8emLQADJ
tkJ+R5LCEdc6UBpVxnFT7rnaOLMm8vXIMXjGzZuFCaQvxhXEPAAt39o2a/uKz4Ud
jJLOYU8h3HAGCC9+8S9JjX0obX532ioacg0lSOZTPHcULBri67Z2OxQcvTP2EZXy
fWT0aVoTlxeNumOb84OOnh5O+tIO2aHdbKw6XAdu7jgKJp+hf6BEg9Z5jwGZuzYJ
uDWrH4JDLsYvPA8QefFkFZ8Ne4wcx6eAk5m14j3i47dBpLIu5fJ8Y2a5VbwYVW9M
B2ryoEmkz+Z8se2RUJoFbvZQAV9+iRLOOrBWmVebhlg/YEZXvcCQDWOKTLjcccSf
hwtvCamwYpQ/+8N9CYAAb8fFdQ43bOPkXjuClmCj5duE5M0jPnciAzck1pMsa6xh
bTahWGGGWgMBVJZYYizmBGhCPJ5HNRzLeS0r58vYdGJoboYLbefIduuttXq/xvlC
rkEccbIDG4cTJgrKKH8nPZNyXhvtKpFPRk2C1bCvHdONxgnCnaFOqoJnhQt7cwUd
/+y2RV9oAhfODvhiNttyhuC/9qNAnxCsTosRFf70OC7YtbDqlwd1wp0qMlluhGrM
lA+wkeqoT1Yuh9zRpr57YUUe9pW6itQTJDYRPLHtMQzOrxJVt+xL03fwuiUA/Gsq
zB4apPetNKRmkcvzRj0AgEFVjFMRgk3GKBwnoqtVAwM0RAPMsE4nxsonjZEepM/L
LRugtz4S2SziGtIdHD7n5JkP5VSdJTDQWXra5UahWtvnZr4GJAaE5ekzZO5PnzEg
cl3HeBjCmJPwTcLvPp0GZNcSTUKtvhIJXFjO0axqoQk6qhCx9ybTRshtk/E1r6wW
4AhN76mnTXWdQ4D3OcZ5SCtYPNLX7l40BrPMQIbUr2pHidXgCsIFUmPPFdTtOsim
4QeICA0tnE6kC4ZTTBrHA/++3XYGyjPa+Y/xMHwX/SM5VbVxbbGIFnB1CguwUEUJ
N+aYfii3UrSEqaT9/kNe2zVbV6ljk4I9JD2oXg2KNVxTTZ+fjOf9ceR87v6U4oCR
dTEjVmj4NphyTQ52Cs/WZUP1LMj8pPUpdW32oxgfukoNRu27fduq9RgafVKNbKxk
Nzwq5nLNEc1Jy/uxdzYDFzewASopq1lVGc6nHfyI59bgWr7/7rF9/XPrGvQ1lKof
WhsPOjxEDrifWyyJXKmzOnErvtfHQg4JpxKbnLAhzjOvnW37jZu28AROPF7sG2NT
ZYMzLo6qM+iEtxUN8MKx9ahdCJ1ZccORlRET8tjMIC38TNERTiXfSNbWOVzQcwYR
mdtOFjLpLcArbm7bnAmlgeFjqJvZtwfbHdJ2cnLPwqEil6iUywl/kfgakbJyXd0D
GAUopz+JT1Dt+DTVXx/PsGaPSf8Ftblcuk4qDpi6Ws2lQJbeGIgCAlmKiArocUtl
OYKFlK6MlYZJ6hulfLokfrYole8XK+PDa0gmOS9rTsfR8t2gK+gSVfclMH1g0xWa
DZKymzqj55wFLN8s9dIw52ZKYvE57iQrUS5TwKNyHN7yZ1xsEUJmz++XZSgTIKxw
T0yyEcYflvZMntPTOXHVnAK+d+JsUMmW8MC8N/+hGi6Lxd0uUZtF82jWyKVX/dqH
GGAyrgKWl1BDZU/h8O1NqvGWE8LT8uf8n4JL0mgszg2DqkTt0hLAMexfCPlXgqhn
dFcyo4CQxzt/MxDnuuG2roo+SglTQNiyMJ/7ZtjaHsz5PKIRoH7KY3U8weSp6o/3
oWhHp0hZqJj5+CDfLJdOV5E0DD3iURJtMJGhBaHyTbZqkGyp6LceQLvFjoNxjXsY
4Ue20aP2HTQ8oJzm6Q5FGxrGeA6zzMwQDKpwvsYF6V6QJgRw1dvw9vYvhmr8aJX6
ng+Jegq+Xh/D2fTxyo4xe6LCsuF8+ZhGBO0JEw0LR2aAARk7oXiYfCx2JIDq4doV
1e31YrDA3kvxQAa9ptLhJuPAJar8zDXrOMh+1OBp42bNZ9/2CQpCqxFQ4nldXid9
rBGbyUPd0RB7ktD1R4B8PjH2FdvnHPothrq3Gr3DxJU50T08ghSLWWgnBLi+gDwj
xnylulBRdnD5aeGpYw74PjOr6FYnBfwr1NObik899bv16+JJZro/oCEcZNyTGDpa
Ptr1C326qqA+ZxlHdalC4Z+txgw6f/Vaf/kppY/pcTt/Ou5U57poXzHOzV4/4WHS
u0Z8pkM9vUtNemwqRysHHjDRjagZDHZmGR/pNCA0uRaFh1WVJFgbOlQFy2VnJQmu
35M2gijVNBtvhtcE93iw8MV7wNC2E8tzqLLzYS1zRj1tLKiXPKnxB8qJFFLyPtBs
Lu9nRVbIWzV5HF2ZaeuYNOC1K5pHk8brT6umpUENQ1gNOSMB7eMGXIIWrAMTyhSa
V7GQffj96fbs/OuHTm2BPMci43Ookv53yxRwt0/Byhgo0ne7jq/JFNZPMt1K7QKi
mSXc+0EZ0MxwBfipwMMJSWt3jJCEK2doNxSPBdPuZt0hvWLT2aqGL8D5oTJo/g81
SBksKFt3Qd9dHgmi9Z1BXMBTLBgxztfq2gotU6fmZ+t0V3gtR0vbrBWwM6vPPq1A
7XODCIbhbKUMtNJJ8oqwPHuwtDy3ZZ7Hu7dKVNbuJSNS/ElIQklFKkkz7Ept+mhE
4r4ZVUnOBo0F2IFhU4kTjuAQdsIfT60RKiRWVddm6a00TbYmnkGfM0Xr9h9RYgyi
oJBT9A8MfDTV7dfVjpO8Bt/2gwbdY7+MVsoYyboWqJSHYNX2V5InqHvQ5oflFedb
B9WzopUjiIWzmgfubL7SGhqTXqt6sNunmw04WfcrhEsVOimPj1bDb4mm/x3MGE6U
x1vBXmI33ITy40OhUxtMrNn6OhvO7WxEk+YNBU/EbEWg6G9FRBwSQirh2LGK2iYT
eObXWK1V7jRE5LnvT37krt5ZMLtW/2lZ1A29Fy0EcVQ5fO1zemKY7wq/APV9KDBg
6eACi/p6sHsVEtGYGH1vEQCLkFPa69H0RxSETJ0KuxNh8lEUhXJDf4xl1FfPPv7J
u5pn8WDKujkVb6U0c21Dox3HYAh5u4t5kZ3ZafRmOKkI/oZ7oZFn9sfFObZkqVyK
dqeTHuiRBBL6fO03LNsTeXhAyIMMvBZ32dLQcn4klFyF9DpkR0h7X4q/G1x7vNE5
mnKiZnjd0Jm6kxrkTp2h15cLpSfRDdITRcJJV5jDkiCw4c5qRh//P49JM54eZX2F
vwprpDsnZScUt5gmcXWqBNg05I74KJ3oNvML3s+AsIPNslaIa/yWf1UU1h7ltash
tHdGmNgCI361iGd/WhPTFzVRld2cAWwP0UwLasy8xKzXEqC333v5kerHhMJxGkk0
IdR4KrJziR4q1mwVLQesEpV+SgpM03UgvHVl8g3CKOzGRVb0F+MtIXRpA03xd/d0
vbL3OAEceY9xeiME0+6FgVUO6VLGTtRrP4D+P0rGWVwcgThxEffOxFogiugaSiTY
Tmm0ATkIpCAdh5P82Hmb4FVUc1Iflbm2YyGxX2+1A4rn3sdZ7KyIlXOStUG3Vrhy
fUKUbTVHgQ37ddFq2YW5tYenrVi7CdlUbSjr5Vd1SNGabynxPig9qcA7CscnhPEW
OxSIxhnr/pLTdKKFDHv5brhy3EIIpVjXiXVy94Rna/zbr8hcC+GtkxkZ95ckoNMl
3hNy5PXyPFnDrdo+sHOrn14vgaUgZugvAvdUHiqCgnWQ3XYY8AzZEvkTZAtaLylb
3ZoZMMrk1Oqi0dHO6g9t3rMGywWbPFLW2I4bBxGHNhRfw1G44FUI4DHTB4Fr4ICs
OmEq3RAWxMobWhOpX47n5bgRmJ5B1Gs3OA+THeWHMaSOqtF15umsoEvZeSGkrlzZ
srP2UGpnOa7FUa0Rc4A5ENdh6HXy3OSjsAryE1moI43KfyLK5RyluyOTmubQVz6i
9XGAg3djDgipWWGOyuVxm2Dsf7hJg3nARX7IY+pXfJAno6uJrk/ePoDIy+my6ZvZ
XngR7o7rcArvjVmTqvHlxGAGgI0FJm3tTpeu9kZarNgRgS3qhVoDaWafY5aYRhqj
yJCzxeaKV2NXRD28lSJC8K7GDR1QQpOedcRT/NQbMWGFycoXOgB0miZbwr5wX/Mu
oKrwD9NLJcvsTP6zDDrbzoRWK37jHxQc3bKaCRka9SJqkK1uIda/hTwfyAcIeH2L
QVdaUshF8nVHFc9mU8lT/R1QbVtn/S4J0OrYmNrI5q2YlcayQ0aIaIYEDxCSd/ZW
tF+T/W11r04s4PxN9gLi8vi4UwW6sE3H9uUDswubiPnHhapBW1ZywTm5JisbSmOV
/aZH5MRGB+2GtdUEFq3NBJwBlfkiJt+okJUbpcghn6kc578OAeN93pJiQ1JGIxXC
C1nC47h5qfJx4B61uFKjsqfaoo2IYQJSSlb0CDqFVmZbRgZlDZYIjAs3JskagkYX
pe3ryNv/HzVTtZlS4zeHgXz0XirNtauO475c9/H1rJ7YbdoV1lVbCSFp95oA0rVw
H09L9yIhn+xng8cA/SAHo7CQSUCmUiBz+VIOeDAF5t/N4/7kl97QCb39Fa8SrZbw
XXCom1gm2vFonF5a50ZRNSNCirtDlc7KcUrcbtq8P2mOSX0MKjZ7PlFDrJeFhGuU
S43S3ApCb0GtKd9FaQjcF8YSG7ty+zabqtxOKw+3EiwShd3v1rTI3vSR85QmYVJl
n+U01e81FOjM5zfrCYSfM9r2yYF9RGox5gEG9OIVNHwmKCWBeu3ASkWqPfmcjgI8
4qZ4ZRyOxt/HdA5b1RoiESNsMJimXhStECCyno6SZDLAVon4JmT3J6xWas88ULsA
hStrYEyzCaRvclc1BzgHQSnhz14ANeBD3pYN0jNowqPAIeq2S2DJFUHfuTg5mtTX
z4R+x4QPdyFKmJhu7gTPMLTHoS+kkSTCuIlxwXDPMAOErleX3/R3Sfy2nNseQBbl
P+rOEV5yOBVxTiL6PGkCx/CdUbPuWEd48LjWGsCaQKDppLbY9mFmWv9k94Wl+y+n
coSoY1x8mn7wNezCx6ZCm1zGiZCHOFlUxfciDu39Jh0aQm4YDVtU+nW5dnUg8kCi
p16bGL9ZzgNCDmFJ5APB+drGxmCcGgwoC4NOvN3o2IQjRx0zpiYqJO+7U6x/U2gU
GPUPL+i/mSkEHJGLqfWiotf4hzHmUEc2qHo4al6e/UeWW1Y5BxI5j/w4+et4iHpK
8vup127ZxuOoUF8GLrXsQiLEWmkbIQEuFJMKCyrsp4Fy6av1URNx6eCtgYCar8wL
E48IsLF4VC7uw5ZjyxNnLkqA1TVD6MpEs/ViWvQyDBX/ajYYBbowVEzTYpMA8Gvj
JDjTG2g903iJrCurUycWCkMNztLuGdkpHxk/0hN0BxqOhFMtUirLTLiV9BrYK17J
BpUXXxoXAIcrs9HhTUQPFeG+ssuf2uu/FVphwoqn5fjlwTB/c6KyqT7i2uOMfdHA
tQ07HJRrRX5UwnSjFUaIMK3/1ctRnw2DgL4VVNWs1KoGINBBBUjt+/Qu9sRAW44d
uz9f4/bpcSpkNp+LA6LN+6dV5gaO4hO9bTcqRjh69yaegfVkMzHYbHH7E53SV8lf
oHB/pqrOTuBrf1KIauEZXbfFk94IdCnptxIcjp01ux+9GtmdSFogJBAFqgyCInSG
Ym4uv3YdtIrYIBaweIDfaBAp14g7Vd+surfsafXHZmVDqdteu1u30IzBPJsDO1Q4
GCyVVLqGhiMYZ9MKdfAlBuOGrATPCdOeeZLq3Tszw8ukHtm9aNSw1Xf9Gu4unzvv
FAZWLVgMf8m/1Td9mhYwjcxTn3w/PUa2c4I5ZA1rgIKfObRcei8OkZXKzFrryqkv
2Xon4ZLbNgiNDhKDozCjECC8nsAhnE31QMmFM2LRNy12xuvFqi1GpLzzWG1Vardx
5vNSmgyXufiPaK7AGGPuKEaX2Mvs8Yr8UV5Py6PYWCHETZn2sHou43ag4r0WKhaS
WWtJ0HRUbEQ4DBjyy0NjAUUDzR0EAEQoQxOvrYYsM2crG988VKZB++F1IDf6AMmY
TJqzxAHn+uaYDJIaYK5VJI4x8IvobpmFfMpCbljhIXq3ECqeVh2ZTuYxp+4vURgi
1vCIgrxG4wUuFpCekODdTjwZT/M3QIpRHUpg+EIWxuKfvndhqTiBWFHn2mLkzByf
2sMH7NoPA3l6ioySI0juLX5p7TZfyYbxqhkvxB3WQYDHsmeo+xuauzMAy9FtbmFz
ocjjZyv0k40sppCYtb5uX5Tsl1N4V30Y4s6qFLJjKJoIhpHXq/rZpXUxjzGowCct
/7+H+RnGhF3aNjMmVe2Vu+6EC2ySx7iKlrYpVri+EWmIhHJ0kbw1ovkv5hh/SYoC
SVYxP9q2Ag/HRmbpnLvbqqJvwSRzD/gE8KsfHtrahuFh3gVKY97Nouxh7ARyZzjY
cmGmRvqoytlfJiOUGbLvEM0zgXAaWVqoRZf/91ImKOPnPkBusosOTsnLvLmyHHnc
6+SZrETdNMLANw0EjprP4W3dr2CnbjsXXPSrvViOEBK/R8iMRcCpYNR4kL2mOOrs
KIFFul/Wd7rCS2F0nYbOAPj9ItRUF5wVZmGMkQRPakOBvI6Jzj2CGdaitm0pQ37L
QSltpsOQUdeqK6AkZztwWjPn7uTJS8H3mya7qV0b2uSWUlERN3dvmd16QIS7OVQC
QnyAitKj/Ltm5/BuYnUIX+lV+AtAcH/OktFIz17jEWTpxYjPJ2KGadPQWKlrQdfD
0sNpDZlYOhhfH9dMgLPG1BSYufyc1ov26Q9RbtCKaAqMZwB6gbstcCSvxAQ0R0zu
W+BeZ5cG3Wf50Iy5NB2oKm4GDKL0/zxXH4IQXmUNGHqTVTm8ohAroMLsiK+GXakk
R5vKP6QtPAmcEzNj//+brVM0o63be0ldya8QJkxSBZ8HoTKj0TEFIFlaNToKI8Qh
vidl0ErFDhg8R7IDkFwsngrARDPQiHaJWwiQx4aBdQ4ERzW73I5my+ofKRaLDfCG
SpWBHe71zyQfPJG8/BFCunCGczY1eGucaYDXhj+VpWUWQyRFHONMx581h5A/IjHR
7BxLhDjuo80FTy4yvXbO6YTGn0mPz7sJMqXYXHgoJE45HkOYPEeTvrfR0qQZsqmV
xmjsEhAUwiJsLdqs3s5ZPRVcl0l/pdmH0ArIJwP8h1ZmyjTS8UlCX4FHwfdEditq
c6xnG8prz/haKmVPRUmXzpbA3aK7atTkSrceJ/DtwnuN/Eq5dgZ2x683SwhSef8H
w9hbIhtIX66D8/ULRJTQCsB6OcO0Ab367w74hQDd3CyMNNn57cf2FQ7EDpUGlMkM
6OWx2+CbdBGnR3bJ5Dk1sLJvoytl6NDy18HoEuQoswMzW+9bvteO3At536pMVejm
etldQbcl0dtA4VjHfBZ1Z8TAALNVnT/k4Hp2PVNmnuJHXefL49Vo3ipt45aYnfOa
yLk7gw0kp9vH6ctW6DtFqZiCUTC3VvqOy84B3WSrhvqC0tlJZkmTxHOxIrOvN7W6
QozzTQBjbvvSkQPx+hiR/vHo2iuUa5PqwD/YeZMCVt3QVLkkEZzWNgbQRpEZQ5Ey
amFiMczkwtnyj7jS2OMM8EDovWREie97Xs4wDaxQp0609bWgHtaNpEYQE2ERWvOE
R1TP+lEOxeKb/p654zNUswgSWeTbPlo9sOzHiaLP1XtbRNnU0OLwDEJvCQxMSUsE
S6EUDB5TXx8OZDgWWCBoAaxQwOjStLaCiHR2Z7ONcCtb3p+UEWFrKhxJ0CGavelO
BUrtYfgdGFAmXq+BH6yvbnNByoEpgsiZ1V/8n54z9fyPXa93hSmIwv5NLppjpxrx
yVvQeFQ3ZTmvXY5aH+WQ6T6C7JZ+yMsLAN1EQxSQxQtQeDAl92uDRrQPiZ6zNsGa
cLGSJz4EBLXPKNQ+FFyZ++uc32LoQOzbXco0cbhHEtb72V1eywPKkTUcGPcAXb3n
LIafm5jgz4BvsKYo0c4Vy1gtP7n84n8Uibvhq+ZteyaKjk/kEnxuDm68fJbVCI/8
vltDBWzKFR+5+Rr1jLetRWTGgroLiDUSLlSwpYGHTAAmOvJX9FL+fJ4OhsUT0RZo
WWjxudoiblz/b/UlKmHRKd+keQe7/vaTxnLfXEzqqaPEq/yNCQtmUvCe4On7aMGu
xHcRmnQ+Gwlr093ll0ftTMEjvkpZhy5YE0vOCb+HuJabOERw0w6SvFVAUWdYwrXz
k6Cua/VEfaM0qR4xgGYeZQ5VV1AyNk9QrxpO2G9Wl6ul2ReAnuKsWP+bqWqTe+xA
xAPFaE5CiMPM6EqZKSnaNZ5LQLmjXLnwws1ZAg74u5uCKnH8vT1MzPuBZSBhugXq
7dvZR80Iq9/XxNleyK3UXPJYhUBg3tHqLVFDtCpFDxlNk4yzRo/zrRvAZIg3asru
fVJrvrhhm9fq5gErw0q/8unqOvCqcBhB5zTX0JxH7mm8/nfd/ghQsJ+T3/0I8WUE
6gLXuECt/cF0PMLn2YipJ+XbqQ1FIpAymgeK4q/xc1PdNdXTs966avsIrad7ARHb
bKqztm6QOcMARojSeHEJg4+a64nxMDAPwOG2YAXJh73LKaWl44A/FN4+4736s6VY
d17kIa2Y63b3Y22ekT3RI7TBegX3fVG+Yo/6SYmERy2BZ8vAwRSPBGBxiUgXyVhY
mqQmMjwe/6TAtY0ATtHTxTUXBP2BaBezQk6SLT1NLFGvjCgkIW6nuOdLeLeBLi9U
fbCRfELJw0ARPdfbmKagPg/ZpyXBvc+ApFpk9lU0h4I34LIdk2Bdd785/ENmPurW
f5Rla8OaElrEptuwpRomCn0ajXlHK74qy/gpgnHdSgJRVUcm6PngtMugWiJ8qUDu
RNVZTURr9NdfsMrvSeF7bw6biRg9/aTAHs0ZkjXqCqDEOC7MNs5/ajhslGMil0sS
8jgk+QuHoND7Z0Y3u8YrKl7+CBiYvHCvh0Fs8n7QfAGHqVoeGetOHWSv6urBshVx
udA6gBI0a8v9zDAggW0kp2MzFlD/7VjtmYGccSkfFTVwFkbhQv0rTxZuoxoF1Ydu
wLl4jfUuPNmlFgua8tGnRSs8Vf68/+Y2+cGK6Hg0hTfcYqLa6bnM0PJu6jv+hUmv
63UnFf/z1rnkgwLm8PnJvo6/hK0VA/79Rq3WTlsXhmPwoPMLRsTeDFJ1GUw0/Utk
WhfqDhRj7+rnDstuAesu+ihlwEV0Z0glaVVsn6FrP0KNIEMEAmoSbbsWU612x5zY
xJdM0OSyBBsHKcjj9mJ2/cACJniX64GyUG12vB5mNa1uwBB6BmyLYBZnw/XT4V3/
S0ePT8Ae+0UUt88fB6KNFwtre25a9HJeO0C2KDE+AchkdupGjkJdy18mO23KHy5E
/e03znwZgZ+MONEEtnI8ZGXLBNIJgj4N7bWSeFby8gHGlVbDmLXA5sP8XsiR1Lba
Jf37gDhl5WrydhCKnlr1DU73Hqqlputv4/X98bd6kLX9gVFcHGuPFWczQaAHoJQV
0orvACKawRsra7POZsPtzP3zuoVWnVrwFUoz2N/T7AjnM4Z2G7XnFVDxirKPj3q9
48gv9CtUhnKrOmW4Mfbbf4Y56B335c1y8LOyf569Ul8a6/oORheUYr8OJhscWNsD
uW4YkBmgXkP3rC/PP9Lxgt8xCLAv1G/eGHUDrZ7sMVomNhtKpphO4MU+LTgFiikf
LXFCHAqBm3NUZgRpv49JzoWAgLyo359UPWfSUK6jC+/wMvQ3FZ+eRHRsjZ0mgfRw
Mz7GmV+OsB4ok59v2cOCVFdmefxRz34JXVefrhfje4uvEBXmIj7iyT7d1XRw8+15
HCqRWpKRjGNmtbrphI9U50oRzDpIvLO59zFTcSW1ZRhIm7qM2ounIrsiHvd2d6pJ
PsGNEea+a+bsrm9Jf2pdhSdcfdq07t0zMJLnZApEn5nHKS+ve4aUfngHeqG3s7cj
YwKhHzdBGQEY6iJiRT+VU87IrxLoFlVwpceCD+RoIHL1ZrhIwH95pXY6MzLVIGfL
Q/lyUmdngR//3FhFdVnMl42JT2jfR5BKZ1bmz2fKZ9BHD/IzlGcnTtMFyVMtAvFP
kOTNBFXqzo3naWqX/qslCujbdpmUQdQoVjgWGgux28U/eUJEzeg08X7nAiDkHOIX
FEQMpkpglbg9NZ+FEFZqgk2PqImiqrL4GnpnT4wA9FZoLFBuTu/vpRD6320XMCpr
cx1iB+d+LyJcf5WSApB1w+UKj8Tvk1g6yyG1+LfuAxODU634yBjDLnJuk808SVz8
Ad9SKNEU+mtCtCTRUkjtgkYr+alhl4s/Fznc2aHxbgUVObEZk3hC83C29w3tsio1
FAfYpocA0hN/UcchMhZxeqVIaPIK0PrAyMFrbJedyLwq/FCtj9qNoKqmX6Gh7pnp
vG9tysmmVE5E6AhaQ1l2/BlWWjNmI0WGupls7xtxWWATslC9H/FcOrxzoEBoBHnO
XdhuR7zWZEgQS5xsjc2fjir+rAFPWQ1HoW639U7c+XbGHRfYach1F/kMW/gfA310
IQjEHuvS0Ro97OLrloY0Byc0G6WLjGF9kUPX1dQPYRGBbD7Zd8NppIOrkZBoL+ss
EceKR+wOc3+CucVU22E3Kf3Crio9+87fQVudv0OJFTR17r/vn8dAji0n05KiOMEA
nymwaAnDVuxcka0yKL+RYOI+J6xOK7TxuWPXwEUTdjHVgsa62QC6P14NuU9MrURi
evgz47HBNiFKtuYT/1STl/r+rPALAGxx1U5OccanUDnOjHsSOXr5hK397ZSE6RBg
kTtnri16sI3r6tWbKbhkfQ6eimWf/IkMDJCdMrpnxBt/RmaVXUmAvk4fS8fPTCEL
FoRNPVbhzMfblxZnOqFsEbzAPiVqChwlNiBenuJHU3WFmMJ/7QWRZoT2P7gGWMtq
XHnXGXVnm/MW8QEnRyDFnZlg1lEIRBRduWGsmCCHr8h/P1dEo/yh7Q4aXI7WIznl
4DNxis0dEWAUPxH8UE9eHfXZxhRuHqCXjnfrj6K7/BTw+thT3UhFKQNENzOVdvUe
nSJh76SPPIfgUH5dfEQnVGfKozZAcqv2CwnjkEl6581RhqEHYfIY++XzzjcOM0QC
aB0Vx68kjxDU6Ma95pPqFVolqrguYgjlNyaIbUmS209wsPX33zbfTz01vr04i0Uz
suCnvz7KyJzLLTUY01B1Q3XvPB+qr3k+R82TPJOx2cs9D04q+9RZsPD3j69AWIEB
wnEg+PfvpZCL8FQ3bgQsM64xV1pCdvXAw0N+1Vd9WfZ2ebgP8HOZ0wL8tZPzzxY6
adE9DmlVP3uM9DZI6yYNNeuzyP09g1XX0VsYVoxMtLQ6t9s0Fxr/YLXRNs2NPUXX
skOjAHNqT1Lc1iir3ltrPR4tdHUf23HsNddPDPmCrGiVseTEkEAV1qv8IJ5tLkLJ
9jDMIQbWdq3qgaUfLv5+u+XVFfPqYHKVBVUfuUYBRV/DT4hjASRmmg3AGh3e3Twd
h23mxwFi3CyHzFM+va7gjC930QUW9g9o1mQE6ezzjPZHEvMRkQqny3H5RzvGDmFK
+r/OaIjFnVsbLf9a8t2LDv91rEFMzUULsBnXKz5i6I2nUdKq0S3mF6sBIgFJLhiw
ZOCffrmHTSMTaW9mgjqvfBpCm+sHhQ2+N5NllnDvK4oAMhm9UZdyYJQHb+khiplX
lQu3cUMlAXtv0215BOgMTZ5fhRQtLyrz3XKEIFYO+HdEw1/jZMCwNT39Z1rZzNJN
6gbhI1fCbNyf+R3IduS2nyv3L7cLDw9hlYdBLNcGCzhcnls0YKu0Pl3XfxWN7xYX
9uf3uOsX5N11G3hZCf2C7p74BgH2Cq7pgNqsnBIxbY5wLVAjXibw/WIEt+3rnb3s
llhQgmVbi99GdAmUHSIGF8gfXzvtWoH+UFGsAPHWZNdg7uBD4nTSqy0Cz6bwSGXj
afeAYdwBMbTWs9w6aE7IIdqIPlzOeunDr1Fgh8VZRwVHpUrP0KCcBBzk/iq5xx0e
0DafvOhJQfgTwzXp1CJ/MyI2glODzL2bVM0dagLhbf+WD+aI7BhWxxsMy2+7Lm8X
W+OXj5Y/bhTmvDgvO+DgPhKsjKdn/QAqNrzTTYQq6J8lfPG7/2Ufpenfs6xJ8fUW
lUP7IiqGjAnpeIvhBaf8ODt0AVfYGVuFZv0f5d5FJoKZ//5hRZyW215d+U2sfOY6
m6mscuFUp+AoF3Qu1fHEbRLOFdxvfJPHSoO/kM1az0f2yIgmoA61Lf8/HFAHThWv
s+1Lm17oqg28l6fXStyxv2LD5sA3/5t6+JrGjpbE9vANIuhfo8d2EhOfD9VHyGzw
HlJhVnJ/Cq2CAxWtFsU3j/n1VSqxFA8nghURassIWe6caamf04gNd0Rl77T32oS/
txILqYYvG8osSEDl033i8LxeqaqmKciQoCwEBk1RiGIS2HlOctcT37rIQtUq2Z0Y
ySdBWGccJUT3OGZYQ75NmXbzTHg+g3EaqiWcPKnyMciovwOd/zE64TPFn/ANu+53
o7sVfNsx6cxFMi+lWbqN9AOjHQqmt+gW69Ffrq4hW3Ew8fNAUiuP+BaRNSp83XDS
N0k79Txemvb5Uth26BTbLwgrny+jKBMi9XdAcxcv+3M23EQsDnBYDsl/VYhYuyV7
m5ivQJbcJ8RWpZxDtI02TFIk4ttvLNPClgyfcQYOrBaDHBUP8BQL3CQAoEUko8gy
J56A5863zLVP5XH29xJdvqmDjprHSWieyLrsOUBAMUiCFV9H3l0kYgqKsuXqjJ+5
63nZ0E53M5sQCNDQxEYq8R0v0O5+yJYQFMQVUSLu30mrpKOSR1voCWq4a3JsFHiR
9NQe2LYTBUbdGQ6mvpJOTudlsjELT8wKKrMWV8/8r21TrOqanSLFPdt00sVLuVQw
DJIMJ9Opp7vz/E0/Bo03SSa8AMzSh7cDNe9tPsLlvvC+OJdi59EOYQ7jGVGYbh6K
hQnZcGcaRGbqAWdoX6s7BEFOom2SBgZ9ba+a9cuzGJr0CAHcq4wnH+0tyFi84cP1
oYhAggM4go7UulSMrnk3IREb1s2MgUp6OhsUybkv3aD+pFCFFQw8DGG+tpVSb9nP
JwGtlSnIuO41R7vsbexyqMYB4brRinx+4/5tHqE5+ujp3uBzdO3UQ8cdKdo9vqsL
sqYEfN4uNixiTaPnggvCOWvUyjKkxurbimGi34saH59ybUmyVc1rcrHjYaNKY0Ab
iTK3JWpg6/1zo1Y0NUilc4zIhtLkS/531rRwQLCFFH0i305PTurApoM/TntvoQIh
zdVS6n+wJd5iHLFxSoD1cFTVk71NdmVoJ9m/IiNp+xWB1N5kccG8cxVe9DHcRjdc
2TydVFCYgVelQNZqfMvtlOC8fGItmtODjW4ETmkH47xJZcl+HAvsavqAGhJwo5zX
rBb/bFwPQD4/oV5abhwre1bF+JvENR0+mA1nAU/qsbQL63bu5e9z8m5PaaP2lb3+
/d6ZW6M1110HVJQwzdldRy5VDQpicFsfNV2Akaa5+pruxsc6/jdR4I/krcD4s7tv
3uNwbgkGLC4WyHpmDh+Yr0g5nm0UKrmfXMm3vSSjOTR+oAZMGGZR21cjgO1dMCEk
dbNtnP4d+3NEjozljuSU1IjiAmewI6ZDbA7NrbhNMGhwnJ9ZZGYILxV+vawzuLYr
eMOTVmETTFE8FX3FIFM8vdxJZ+afEtqCcj5hChHMe25262C2XtNIepZ9xcK9jZs9
61iVnjsJIfyV5FK/Ud8qpj0herp8YHQxQcTPtBel1DiRVWbJfTnMhrNVbK66YmgO
8m7ipoHhfSRjnYlwJyfP3ENM/lwpBblClSYj5gLnOtMvv8UiVOgNwFQhlGvbuPw3
+c2JruregQQVGv3KSNkL+FmQ+771aH8T4R3Px29H8vfW4zF/YIgZPmzNRitwK5GX
fRV0cQ34I0phsV0ylMWFbQPlAE7gyN5IY2C1q6K/Xp4oHCskDzgR5YGLVSA8Tfc4
5TuS59PsbL2qu+fddYNXA7IJ9A8vh6eaR2eg0gYISyhTVHNBkZ8SRTjrGxrONBHN
akdB3lB/ywwVERKopC+CzT/3zUmO8Jq0sBGowfUv8qvAXa9bkGspsOEXACWrZ3KP
7giJy7miZ7MKq3g2IZzJBTNlbmmG9OAho6iUMA33xqw7yeNwbbjk8KLCdQQ5E1oP
EoaWtEu1Smw6FDg26tDCNOnRGcoi2E/g06e3vOMWVIXRYzTp+AudSEu0DzeV+zC1
KM3hXAK2RLj1Oh7yKfXxNsFqmOOBm7UREGBtQlwQu5CHcaU5Ny9ytyZ5+UUJ0a4N
FUUG54I+lyVqZsXKlIANQbuId5QCNGT5X80MGoLIdZrY1wwDVv9qRZlV1g7glyLP
opPfBRwYmzsz4xbIBLzBQrHK+NDOTQzaifaB3MlNhwiBTe2E/7iAreEXXzaX4s5f
luhJwq2eutfB1sU+rC4hFCparmPTVzBmdsPe4PogwjGngL/Rx+YkWyn+yp/Hk9tQ
kYysdgcX3OlX1TOn47L23F6EhxSr7AVirlAK9MOCFZOkBBcbz20ysLgrgO8Nbm6K
OjvvaVGN1FAoctvfpWOUfCr/Mxn5yIy45wvOLSOiwqiNFiWzjDQdU26QK1OrxEnR
KhuD9TkSUq69145bqbgNW9tgjKEy2kmm9G8h4j9/i5Gj5oQdX7Li9qF5qyNLgPe9
5kJZ4Z9s7unHJvFgLWpwkbcbfYSC7h7PhltIrV3o82nNMMz8aYNA0u1U4dm0kACC
7g7w1RGOrNvObArXV8cQPwn7wYXRndL4/WTZVEypT2UR0BRTpj+PSNH8vmoppHE1
E5MemfDSAKFO3w8lk5ClblmtFbuqkxU5M3CQmGhL12kVbWnGjdvDvE9kpSE0Dyuu
+SkhFmt8uExWBKCEzajRhPGZCz/zBtRDmHxABVgR3lvSRY1R+R94bO83QChF04C2
KKUEEtTqdA6kIm0S67BCd131fGisY4XMXtg4JCu+/eCOp4dP0Pc9j2jD0uYw1jPh
PhFUBpQ3o64bVgii0pwNKS9DujRoUyyMxFMorY4xZIBocKdp/pK0tqx/c0pveQaf
UcubEjT3hBBAxj5XF4vIT6hIebR6kOQd/jpxUhn67AiZpj1C4BHUfhkxuKgpvaPQ
SU9z+8463EFMF9IKkNaReHNS273eku5vLccC/IVdM8IfHxr5wHUbZy7/j4A0HOwH
+tOyQq2QdtEpDXet2PPtmvetbb4oclCsqKqATh+HGjesfu13WqV4bs3N7jMylye3
o0wynjqAbffNCU6eTN4G1mkswy9JzvGzeNQwRoDdbhMmS67bSJ5Zb93DakyWaRtF
XzsskpQa7DKrxa8DvE/b+6nlTRCqRdx5FiNwkaddAYIJXQuDZRACdMBkAkUq45e1
U3dLfFgygIlDUNTV2x0S6BJPII8AK4ke8atlNpqab1ZdyhuBz1LiBVOBVOpJ/6fx
t7AoKaFrPS/TjJriC/fWN7oPCvzqTkSEqrtM2j4QnqeUlBvWdojl8HF0tp4AnGcu
rgCBbrgnsLtxz4Ox91UuI1msofIXRv7ZVy8MQkxsOmer+B3rwdeqw5TQpeLbitJA
AvhIRfrC8R0w84aXrA97DEPIO0Zu97aXQGT5LEzyY/Wh6aULsvFh3n1X+SFpiXfa
VCDVOl5vkHKUq0FOQ0Db9YxA6WbuLKyjCF5z25liq7qAby/KjTJ5eqYcwe2diEBs
FGq4ALFLzOP2WKSoSMZh/MLR4c9aQojfdps2yP4Yq7ysVRR5CYvcfTw/QesrG19j
LQEpRJJFF8I8BrNLnNVjKDAjDNdzYYyrplePINDV7CKb3LmZZ+EtPMs5NYNZmQHz
sith01jmX0eJKFb3jYP9xrZK6QHSLnLJy+L70SAZngppGiLzZuQ2Kp7e/V8PJbK2
+mPSgL7KB1teqKbwuexC4uC9v6HNmgH8zlrFcF1sxZQu7FR61fxfAQIV3+mC6UG6
inrDx3UvcBk0YZWFiBSC6QRRNDvWud400Yxz+CeQQiOhwSBTPTw13WS985whzaA3
Ch6RpzkusM5+vSe2gmOi0QljC7dYJOMJDH+QmvlR3pUkwxn761muPzzmbpV8QJxu
YTIjVCbLAnyWiVeYA6WrtuYVRQ4Q3xX1oLuGqsQiAwGy/THPCC9atBN+5oXNjFJm
FXP9h3GHADGU/DBG+Hj6erXmrUfz831CdNILZrHr2dVoLowNj///XzsvfZuQ2S7K
ziYDfUU3C16OrPwDjLtSsvd6Sez0tODI1Y8Ub6p7XBTqZALnvWQUiYlqMOa7SHV5
BsLuxDr/NjmfpmLAePOdk3i4K9sYec+mcdvam3wHpw8+Xedl+kRJWcYE77v7+v7q
RjCaLx6QwoX4WbTglqwbSRyx2bc2Ox7u9vnxaYQmgm+AewG19LNiIsQbXlOo05K7
haSl2LXFeT9BfYdkZ4hmG5gLImFVZjS+h3qPCJ4jasBSsugKZSnhOkyVV9TDX4ky
RtWnIQGQFzwC539NbUSsIwkiC8hzKpXN76cE2szwBjzRxJCr+9U2I4sq17NhLwMx
85wup+Q3gcAGr4cBEY9VpfQwH6f7cQTulp5vwf1snSDrOoirZXuZR6BJt4WgyCRx
I8hph+ofNhyB3Mm64dYQzly81UCFbazx0PIGeJEvTTeF03aQXDd53iRok3fr3lLd
ADoCQ4p+xXbVfwEjk3i5u3sa6pIkLAO5A0EKZTZaQqu2F2x3ok8Wg+BH95XxHsfj
P7xyZTbtI/Hzv1Tx4y4zVPiyNLeb/Z+YdMeAvXlXKXOor6L/d9np8lJBG5Up7LRi
VMrEYnjUYcZzZntt9j7fHEyufc+bAe/AeXUDGLLiguqJcqq4szKYNkO19scXgaYy
zvlYGevvzHUnch99KUbCgbZxAEFVHoka4ULDNSf/qPadU4m75Y6LWB52UtUnpahY
8Xho6mkrvfERE+QHH0vAx07YBHR3YjnzQ1yHLOPs60TkCqICPYlRRKtQ6CqT1sqJ
d/O2OwzO/fveLfvvTaURitHi0qZblzAXVQlVRN4vD+7lfJSXh6aD8njGogBFcZY5
T6luFL0ikMWh02v/khJVO0A4fzKNAzo5I8RI2tM7v9oeBKX379nNSHZoCiAZy3Je
f7IeEgwYjkO4qeu28Ii4ID6iOwoosf5R6FE0/3NPqKlfu/AF1CH6Zk+mJE1Bq680
ECcjiovv5KPdo6jVNpz1bnmzdY7iMVQtnPzs3ybbb6ixf24eoQkGDSZmBox5LEXL
5b6/WFILy92HCJ8ftbqT8esmvLp/cMkkRzepSNQhnexF1YxYI8IHemoZaRDLeXWf
rO6P64YqCIV2l576DrnibCeOJqIP2G/NBBofdGRseEIfKwzOQe4VrwD/P2gN8SnQ
O2KJwz3W+Cg706BKgp4q1KuwugW0v0I8BBPR5TAFkdf+H1kFkmlZoDnC7zCtXHPp
pw7OVcn2CsJBoJycvOiRr55xgRN0sasN3BP4ADo4ES27AL3LEZs56AFFnJRtW1RD
bO11iJBozzYKeFfPwpxQlSSlMwXMoQXBF6ojP4AzJUZM0NVsWqJxPC8pQDC32QEM
e0VVcCtLZYvCxNpfjPyDYTjiBmFw04EECB2LjNgyZPSL2NEFYRj9LhgTeSNsG2Ga
KvxMALs308+DWiXpNquFpji/8AFfMloz8cbGPl//H+hd2PIiGX7ztnpwi24kDtTg
7RuoYOXWIVP6HSbCsOdqh3rHLtWHd/A6Mox9eWfd9p244ND8BK6MKIA2L5ndeP8P
VPcgNWmCSCnIXw2qROf7GaJOgD7fARJmSElvLqay+3QPEYDUDB4zdP0a4LHxoEK2
JabGSWBBpuFVAJhuxA72rQ==
`pragma protect end_protected
