`define ADDR_SYSC_RSTR                 7'h0
`define SYSC_RSTR_TRIG_OFFSET 0
`define SYSC_RSTR_TRIG 32'h0fffffff
`define SYSC_RSTR_RST_OFFSET 28
`define SYSC_RSTR_RST 32'h10000000
`define ADDR_SYSC_GPSR                 7'h4
`define SYSC_GPSR_LED_STAT_OFFSET 0
`define SYSC_GPSR_LED_STAT 32'h00000001
`define SYSC_GPSR_LED_LINK_OFFSET 1
`define SYSC_GPSR_LED_LINK 32'h00000002
`define SYSC_GPSR_FMC_SCL_OFFSET 2
`define SYSC_GPSR_FMC_SCL 32'h00000004
`define SYSC_GPSR_FMC_SDA_OFFSET 3
`define SYSC_GPSR_FMC_SDA 32'h00000008
`define SYSC_GPSR_NET_RST_OFFSET 4
`define SYSC_GPSR_NET_RST 32'h00000010
`define SYSC_GPSR_BTN1_OFFSET 5
`define SYSC_GPSR_BTN1 32'h00000020
`define SYSC_GPSR_BTN2_OFFSET 6
`define SYSC_GPSR_BTN2 32'h00000040
`define SYSC_GPSR_SFP_DET_OFFSET 7
`define SYSC_GPSR_SFP_DET 32'h00000080
`define SYSC_GPSR_SFP_SCL_OFFSET 8
`define SYSC_GPSR_SFP_SCL 32'h00000100
`define SYSC_GPSR_SFP_SDA_OFFSET 9
`define SYSC_GPSR_SFP_SDA 32'h00000200
`define SYSC_GPSR_SPI_SCLK_OFFSET 10
`define SYSC_GPSR_SPI_SCLK 32'h00000400
`define SYSC_GPSR_SPI_NCS_OFFSET 11
`define SYSC_GPSR_SPI_NCS 32'h00000800
`define SYSC_GPSR_SPI_MOSI_OFFSET 12
`define SYSC_GPSR_SPI_MOSI 32'h00001000
`define SYSC_GPSR_SPI_MISO_OFFSET 13
`define SYSC_GPSR_SPI_MISO 32'h00002000
`define SYSC_GPSR_DP_LED_STAT_OFFSET 14
`define SYSC_GPSR_DP_LED_STAT 32'h00004000
`define SYSC_GPSR_DP_LED_LINK_OFFSET 15
`define SYSC_GPSR_DP_LED_LINK 32'h00008000
`define SYSC_GPSR_DP_SFP_DET_OFFSET 16
`define SYSC_GPSR_DP_SFP_DET 32'h00010000
`define SYSC_GPSR_DP_SFP_SCL_OFFSET 17
`define SYSC_GPSR_DP_SFP_SCL 32'h00020000
`define SYSC_GPSR_DP_SFP_SDA_OFFSET 18
`define SYSC_GPSR_DP_SFP_SDA 32'h00040000
`define SYSC_GPSR_MINIC_RST_OFFSET 19
`define SYSC_GPSR_MINIC_RST 32'h00080000
`define SYSC_GPSR_MINIC_DP_RST_OFFSET 20
`define SYSC_GPSR_MINIC_DP_RST 32'h00100000
`define ADDR_SYSC_GPCR                 7'h8
`define SYSC_GPCR_LED_STAT_OFFSET 0
`define SYSC_GPCR_LED_STAT 32'h00000001
`define SYSC_GPCR_LED_LINK_OFFSET 1
`define SYSC_GPCR_LED_LINK 32'h00000002
`define SYSC_GPCR_FMC_SCL_OFFSET 2
`define SYSC_GPCR_FMC_SCL 32'h00000004
`define SYSC_GPCR_FMC_SDA_OFFSET 3
`define SYSC_GPCR_FMC_SDA 32'h00000008
`define SYSC_GPCR_SFP_SCL_OFFSET 8
`define SYSC_GPCR_SFP_SCL 32'h00000100
`define SYSC_GPCR_SFP_SDA_OFFSET 9
`define SYSC_GPCR_SFP_SDA 32'h00000200
`define SYSC_GPCR_SPI_SCLK_OFFSET 10
`define SYSC_GPCR_SPI_SCLK 32'h00000400
`define SYSC_GPCR_SPI_CS_OFFSET 11
`define SYSC_GPCR_SPI_CS 32'h00000800
`define SYSC_GPCR_SPI_MOSI_OFFSET 12
`define SYSC_GPCR_SPI_MOSI 32'h00001000
`define SYSC_GPCR_DP_LED_STAT_OFFSET 14
`define SYSC_GPCR_DP_LED_STAT 32'h00004000
`define SYSC_GPCR_DP_LED_LINK_OFFSET 15
`define SYSC_GPCR_DP_LED_LINK 32'h00008000
`define SYSC_GPCR_DP_SFP_SCL_OFFSET 17
`define SYSC_GPCR_DP_SFP_SCL 32'h00020000
`define SYSC_GPCR_DP_SFP_SDA_OFFSET 18
`define SYSC_GPCR_DP_SFP_SDA 32'h00040000
`define ADDR_SYSC_HWFR                 7'hc
`define SYSC_HWFR_MEMSIZE_OFFSET 0
`define SYSC_HWFR_MEMSIZE 32'h0000000f
`define SYSC_HWFR_STORAGE_TYPE_OFFSET 8
`define SYSC_HWFR_STORAGE_TYPE 32'h00000300
`define SYSC_HWFR_STORAGE_SEC_OFFSET 16
`define SYSC_HWFR_STORAGE_SEC 32'hffff0000
`define ADDR_SYSC_HWIR                 7'h10
`define SYSC_HWIR_NAME_OFFSET 0
`define SYSC_HWIR_NAME 32'hffffffff
`define ADDR_SYSC_SDBFS                7'h14
`define SYSC_SDBFS_BADDR_OFFSET 0
`define SYSC_SDBFS_BADDR 32'hffffffff
`define ADDR_SYSC_TCR                  7'h18
`define SYSC_TCR_TDIV_OFFSET 0
`define SYSC_TCR_TDIV 32'h00000fff
`define SYSC_TCR_ENABLE_OFFSET 31
`define SYSC_TCR_ENABLE 32'h80000000
`define ADDR_SYSC_TVR                  7'h1c
`define ADDR_SYSC_DIAG_INFO            7'h20
`define SYSC_DIAG_INFO_VER_OFFSET 0
`define SYSC_DIAG_INFO_VER 32'h0000ffff
`define SYSC_DIAG_INFO_ID_OFFSET 16
`define SYSC_DIAG_INFO_ID 32'hffff0000
`define ADDR_SYSC_DIAG_NW              7'h24
`define SYSC_DIAG_NW_RW_OFFSET 0
`define SYSC_DIAG_NW_RW 32'h0000ffff
`define SYSC_DIAG_NW_RO_OFFSET 16
`define SYSC_DIAG_NW_RO 32'hffff0000
`define ADDR_SYSC_DIAG_CR              7'h28
`define SYSC_DIAG_CR_ADR_OFFSET 0
`define SYSC_DIAG_CR_ADR 32'h0000ffff
`define SYSC_DIAG_CR_RW_OFFSET 31
`define SYSC_DIAG_CR_RW 32'h80000000
`define ADDR_SYSC_DIAG_DAT             7'h2c
`define ADDR_SYSC_WDIAG_CTRL           7'h30
`define SYSC_WDIAG_CTRL_DATA_VALID_OFFSET 0
`define SYSC_WDIAG_CTRL_DATA_VALID 32'h00000001
`define SYSC_WDIAG_CTRL_DATA_SNAPSHOT_OFFSET 8
`define SYSC_WDIAG_CTRL_DATA_SNAPSHOT 32'h00000100
`define ADDR_SYSC_WDIAG_SSTAT          7'h34
`define SYSC_WDIAG_SSTAT_WR_MODE_OFFSET 0
`define SYSC_WDIAG_SSTAT_WR_MODE 32'h00000001
`define SYSC_WDIAG_SSTAT_SERVOSTATE_OFFSET 8
`define SYSC_WDIAG_SSTAT_SERVOSTATE 32'h00000f00
`define ADDR_SYSC_WDIAG_PSTAT          7'h38
`define SYSC_WDIAG_PSTAT_LINK_OFFSET 0
`define SYSC_WDIAG_PSTAT_LINK 32'h00000001
`define SYSC_WDIAG_PSTAT_LOCKED_OFFSET 1
`define SYSC_WDIAG_PSTAT_LOCKED 32'h00000002
`define ADDR_SYSC_WDIAG_PTPSTAT        7'h3c
`define SYSC_WDIAG_PTPSTAT_PTPSTATE_OFFSET 0
`define SYSC_WDIAG_PTPSTAT_PTPSTATE 32'h000000ff
`define ADDR_SYSC_WDIAG_ASTAT          7'h40
`define SYSC_WDIAG_ASTAT_AUX_OFFSET 0
`define SYSC_WDIAG_ASTAT_AUX 32'h000000ff
`define ADDR_SYSC_WDIAG_TXFCNT         7'h44
`define ADDR_SYSC_WDIAG_RXFCNT         7'h48
`define ADDR_SYSC_WDIAG_SEC_MSB        7'h4c
`define ADDR_SYSC_WDIAG_SEC_LSB        7'h50
`define ADDR_SYSC_WDIAG_NS             7'h54
`define ADDR_SYSC_WDIAG_MU_MSB         7'h58
`define ADDR_SYSC_WDIAG_MU_LSB         7'h5c
`define ADDR_SYSC_WDIAG_DMS_MSB        7'h60
`define ADDR_SYSC_WDIAG_DMS_LSB        7'h64
`define ADDR_SYSC_WDIAG_ASYM           7'h68
`define ADDR_SYSC_WDIAG_CKO            7'h6c
`define ADDR_SYSC_WDIAG_SETP           7'h70
`define ADDR_SYSC_WDIAG_UCNT           7'h74
`define ADDR_SYSC_WDIAG_TEMP           7'h78
